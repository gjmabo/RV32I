`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module IntXbar(
  input   io_in_0_0,
  input   io_in_0_1,
  output  io_out_0_0,
  output  io_out_0_1
);
  assign io_out_0_0 = io_in_0_0;
  assign io_out_0_1 = io_in_0_1;
endmodule
module TLXbar(
  input         clock,
  input         reset,
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [2:0]  io_in_1_a_bits_param,
  input  [3:0]  io_in_1_a_bits_size,
  input  [3:0]  io_in_1_a_bits_source,
  input  [31:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [3:0]  io_in_1_d_bits_size,
  output [3:0]  io_in_1_d_bits_source,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input         io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output        io_in_0_d_bits_source,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_2_a_ready,
  output        io_out_2_a_valid,
  output [2:0]  io_out_2_a_bits_opcode,
  output [3:0]  io_out_2_a_bits_size,
  output [4:0]  io_out_2_a_bits_source,
  output        io_out_2_d_ready,
  input         io_out_2_d_valid,
  input  [2:0]  io_out_2_d_bits_opcode,
  input  [1:0]  io_out_2_d_bits_param,
  input  [3:0]  io_out_2_d_bits_size,
  input  [4:0]  io_out_2_d_bits_source,
  input         io_out_2_d_bits_sink,
  input  [31:0] io_out_2_d_bits_data,
  input         io_out_2_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [3:0]  io_out_1_a_bits_size,
  output [4:0]  io_out_1_a_bits_source,
  output [30:0] io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [3:0]  io_out_1_d_bits_size,
  input  [4:0]  io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [31:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire [4:0] in_1_a_bits_source;
  wire [4:0] _GEN_5;
  wire [4:0] _T_494;
  wire  _T_495;
  wire [3:0] _T_504;
  wire [3:0] out_0_d_bits_size;
  wire [31:0] _T_908;
  wire [32:0] _T_909;
  wire [32:0] _T_911;
  wire [32:0] _T_912;
  wire  _T_914;
  wire [31:0] _T_916;
  wire [32:0] _T_917;
  wire [32:0] _T_919;
  wire [32:0] _T_920;
  wire  _T_922;
  wire [32:0] _T_925;
  wire [32:0] _T_927;
  wire [32:0] _T_928;
  wire  _T_930;
  wire [31:0] _T_932;
  wire [32:0] _T_933;
  wire [32:0] _T_935;
  wire [32:0] _T_936;
  wire  _T_938;
  wire [31:0] _T_940;
  wire [32:0] _T_941;
  wire [32:0] _T_943;
  wire [32:0] _T_944;
  wire  _T_946;
  wire  _T_947;
  wire  _T_948;
  wire  _T_949;
  wire  _T_950;
  wire [31:0] _T_952;
  wire [32:0] _T_953;
  wire [32:0] _T_955;
  wire [32:0] _T_956;
  wire  _T_958;
  wire [31:0] _T_960;
  wire [32:0] _T_961;
  wire [32:0] _T_963;
  wire [32:0] _T_964;
  wire  _T_966;
  wire [31:0] _T_976;
  wire [32:0] _T_977;
  wire [32:0] _T_979;
  wire [32:0] _T_980;
  wire  _T_982;
  wire [31:0] _T_984;
  wire [32:0] _T_985;
  wire [32:0] _T_987;
  wire [32:0] _T_988;
  wire  _T_990;
  wire [32:0] _T_993;
  wire [32:0] _T_995;
  wire [32:0] _T_996;
  wire  _T_998;
  wire [31:0] _T_1000;
  wire [32:0] _T_1001;
  wire [32:0] _T_1003;
  wire [32:0] _T_1004;
  wire  _T_1006;
  wire [31:0] _T_1008;
  wire [32:0] _T_1009;
  wire [32:0] _T_1011;
  wire [32:0] _T_1012;
  wire  _T_1014;
  wire  _T_1015;
  wire  _T_1016;
  wire  _T_1017;
  wire  _T_1018;
  wire [31:0] _T_1020;
  wire [32:0] _T_1021;
  wire [32:0] _T_1023;
  wire [32:0] _T_1024;
  wire  _T_1026;
  wire [31:0] _T_1028;
  wire [32:0] _T_1029;
  wire [32:0] _T_1031;
  wire [32:0] _T_1032;
  wire  _T_1034;
  wire [3:0] _T_1576;
  wire  _T_1578;
  wire  _T_1588;
  wire  _T_1590;
  wire [3:0] _T_1607;
  wire  _T_1609;
  wire  _T_1619;
  wire  _T_1621;
  wire [3:0] _T_1638;
  wire  _T_1640;
  wire  _T_1650;
  wire  _T_1652;
  wire [26:0] _T_1894;
  wire [11:0] _T_1895;
  wire [11:0] _T_1896;
  wire [9:0] _T_1897;
  wire  _T_1898;
  wire  _T_1900;
  wire [9:0] _T_1902;
  wire [26:0] _T_1905;
  wire [11:0] _T_1906;
  wire [11:0] _T_1907;
  wire [9:0] _T_1908;
  wire  _T_1909;
  wire  _T_1911;
  wire [9:0] _T_1913;
  wire [20:0] _T_1991;
  wire [5:0] _T_1992;
  wire [5:0] _T_1993;
  wire [3:0] _T_1994;
  wire  _T_1995;
  wire [3:0] _T_1997;
  wire [22:0] _T_2000;
  wire [7:0] _T_2001;
  wire [7:0] _T_2002;
  wire [5:0] _T_2003;
  wire  _T_2004;
  wire [5:0] _T_2006;
  wire [26:0] _T_2009;
  wire [11:0] _T_2010;
  wire [11:0] _T_2011;
  wire [9:0] _T_2012;
  wire  _T_2013;
  wire [9:0] _T_2015;
  wire [9:0] beatsDO_0;
  wire [9:0] beatsDO_1;
  wire  _T_2075;
  wire  _T_2076;
  wire  _T_2077;
  wire  _T_2080;
  wire  _T_2082;
  wire  _T_2084;
  wire  _T_2085;
  wire  _T_2086;
  wire  _T_2133;
  wire  _T_2134;
  wire  _T_2135;
  wire  _T_2138;
  wire  _T_2140;
  wire  _T_2142;
  wire  _T_2143;
  wire  _T_2144;
  wire  _T_2429;
  wire  _T_2430;
  wire  _T_2433;
  wire  _T_2435;
  wire  _T_2436;
  wire  _T_2473;
  wire  _T_2474;
  wire  _T_2477;
  wire  _T_2479;
  wire  _T_2480;
  wire  _T_2517;
  wire  _T_2518;
  wire  _T_2521;
  wire  _T_2523;
  wire  _T_2524;
  reg [9:0] _T_2645;
  reg [31:0] _RAND_0;
  wire  _T_2647;
  wire  _T_2648;
  wire [1:0] _T_2649;
  wire  _T_2651;
  wire  _T_2652;
  wire  _T_2654;
  reg [1:0] _T_2658;
  reg [31:0] _RAND_1;
  wire [1:0] _T_2659;
  wire [1:0] _T_2660;
  wire [3:0] _T_2661;
  wire [2:0] _T_2662;
  wire [3:0] _GEN_6;
  wire [3:0] _T_2663;
  wire [2:0] _T_2665;
  wire [3:0] _GEN_7;
  wire [3:0] _T_2666;
  wire [3:0] _GEN_8;
  wire [3:0] _T_2667;
  wire [1:0] _T_2668;
  wire [1:0] _T_2669;
  wire [1:0] _T_2670;
  wire [1:0] _T_2671;
  wire  _T_2673;
  wire  _T_2674;
  wire [1:0] _T_2675;
  wire [2:0] _GEN_9;
  wire [2:0] _T_2676;
  wire [1:0] _T_2677;
  wire [1:0] _T_2678;
  wire [1:0] _GEN_0;
  wire  _T_2681;
  wire  _T_2682;
  wire  _T_2690;
  wire  _T_2691;
  wire  _T_2701;
  wire  _T_2705;
  wire  _T_2710;
  wire  _T_2711;
  wire  _T_2713;
  wire  _T_2715;
  wire  _T_2716;
  wire  _T_2718;
  wire  _T_2720;
  wire  _T_2721;
  wire  _T_2723;
  wire [9:0] _T_2725;
  wire [9:0] _T_2727;
  wire [9:0] _T_2728;
  wire  _T_2729;
  wire [9:0] _GEN_10;
  wire [10:0] _T_2730;
  wire [10:0] _T_2731;
  wire [9:0] _T_2732;
  wire [9:0] _T_2733;
  reg  _T_2751_0;
  reg [31:0] _RAND_2;
  reg  _T_2751_1;
  reg [31:0] _RAND_3;
  wire  _T_2762_0;
  wire  _T_2762_1;
  wire  _T_2770_0;
  wire  _T_2770_1;
  wire  _T_2778;
  wire  _T_2779;
  wire  _T_2783;
  wire  _T_2785;
  wire  _T_2786;
  wire  _T_2789;
  wire [35:0] _T_2791;
  wire [67:0] _T_2792;
  wire [8:0] _T_2793;
  wire [5:0] _T_2794;
  wire [14:0] _T_2795;
  wire [82:0] _T_2796;
  wire [82:0] _T_2798;
  wire [35:0] _T_2799;
  wire [67:0] _T_2800;
  wire [8:0] _T_2801;
  wire [5:0] _T_2802;
  wire [14:0] _T_2803;
  wire [82:0] _T_2804;
  wire [82:0] _T_2806;
  wire [82:0] _T_2807;
  wire [31:0] _T_2812;
  wire [3:0] _T_2813;
  wire [31:0] _T_2814;
  wire [4:0] _T_2815;
  wire [3:0] _T_2816;
  wire [2:0] _T_2817;
  wire [2:0] _T_2818;
  reg [9:0] _T_2823;
  reg [31:0] _RAND_4;
  wire  _T_2825;
  wire  _T_2826;
  wire [1:0] _T_2827;
  wire  _T_2829;
  wire  _T_2830;
  wire  _T_2832;
  reg [1:0] _T_2836;
  reg [31:0] _RAND_5;
  wire [1:0] _T_2837;
  wire [1:0] _T_2838;
  wire [3:0] _T_2839;
  wire [2:0] _T_2840;
  wire [3:0] _GEN_11;
  wire [3:0] _T_2841;
  wire [2:0] _T_2843;
  wire [3:0] _GEN_12;
  wire [3:0] _T_2844;
  wire [3:0] _GEN_13;
  wire [3:0] _T_2845;
  wire [1:0] _T_2846;
  wire [1:0] _T_2847;
  wire [1:0] _T_2848;
  wire [1:0] _T_2849;
  wire  _T_2851;
  wire  _T_2852;
  wire [1:0] _T_2853;
  wire [2:0] _GEN_14;
  wire [2:0] _T_2854;
  wire [1:0] _T_2855;
  wire [1:0] _T_2856;
  wire [1:0] _GEN_1;
  wire  _T_2859;
  wire  _T_2860;
  wire  _T_2868;
  wire  _T_2869;
  wire  _T_2879;
  wire  _T_2883;
  wire  _T_2888;
  wire  _T_2889;
  wire  _T_2891;
  wire  _T_2893;
  wire  _T_2894;
  wire  _T_2896;
  wire  _T_2898;
  wire  _T_2899;
  wire  _T_2901;
  wire [9:0] _T_2903;
  wire [9:0] _T_2905;
  wire [9:0] _T_2906;
  wire  _T_2907;
  wire [9:0] _GEN_15;
  wire [10:0] _T_2908;
  wire [10:0] _T_2909;
  wire [9:0] _T_2910;
  wire [9:0] _T_2911;
  reg  _T_2929_0;
  reg [31:0] _RAND_6;
  reg  _T_2929_1;
  reg [31:0] _RAND_7;
  wire  _T_2940_0;
  wire  _T_2940_1;
  wire  _T_2948_0;
  wire  _T_2948_1;
  wire  _T_2956;
  wire  _T_2957;
  wire  _T_2961;
  wire  _T_2963;
  wire  _T_2964;
  wire  _T_2967;
  wire [82:0] _T_2976;
  wire [82:0] _T_2984;
  wire [82:0] _T_2985;
  wire [31:0] _T_2990;
  wire [3:0] _T_2991;
  wire [31:0] _T_2992;
  wire [4:0] _T_2993;
  wire [3:0] _T_2994;
  wire [2:0] _T_2996;
  reg [9:0] _T_3001;
  reg [31:0] _RAND_8;
  wire  _T_3003;
  wire  _T_3004;
  wire [1:0] _T_3005;
  wire  _T_3007;
  wire  _T_3008;
  wire  _T_3010;
  reg [1:0] _T_3014;
  reg [31:0] _RAND_9;
  wire [1:0] _T_3015;
  wire [1:0] _T_3016;
  wire [3:0] _T_3017;
  wire [2:0] _T_3018;
  wire [3:0] _GEN_16;
  wire [3:0] _T_3019;
  wire [2:0] _T_3021;
  wire [3:0] _GEN_17;
  wire [3:0] _T_3022;
  wire [3:0] _GEN_18;
  wire [3:0] _T_3023;
  wire [1:0] _T_3024;
  wire [1:0] _T_3025;
  wire [1:0] _T_3026;
  wire [1:0] _T_3027;
  wire  _T_3029;
  wire  _T_3030;
  wire [1:0] _T_3031;
  wire [2:0] _GEN_19;
  wire [2:0] _T_3032;
  wire [1:0] _T_3033;
  wire [1:0] _T_3034;
  wire [1:0] _GEN_2;
  wire  _T_3037;
  wire  _T_3038;
  wire  _T_3046;
  wire  _T_3047;
  wire  _T_3057;
  wire  _T_3061;
  wire  _T_3066;
  wire  _T_3067;
  wire  _T_3069;
  wire  _T_3071;
  wire  _T_3072;
  wire  _T_3074;
  wire  _T_3076;
  wire  _T_3077;
  wire  _T_3079;
  wire [9:0] _T_3081;
  wire [9:0] _T_3083;
  wire [9:0] _T_3084;
  wire  _T_3085;
  wire [9:0] _GEN_20;
  wire [10:0] _T_3086;
  wire [10:0] _T_3087;
  wire [9:0] _T_3088;
  wire [9:0] _T_3089;
  reg  _T_3107_0;
  reg [31:0] _RAND_10;
  reg  _T_3107_1;
  reg [31:0] _RAND_11;
  wire  _T_3118_0;
  wire  _T_3118_1;
  wire  _T_3126_0;
  wire  _T_3126_1;
  wire  _T_3134;
  wire  _T_3135;
  wire  _T_3139;
  wire  _T_3141;
  wire  _T_3142;
  wire  _T_3145;
  wire [82:0] _T_3154;
  wire [82:0] _T_3162;
  wire [82:0] _T_3163;
  wire [4:0] _T_3171;
  wire [3:0] _T_3172;
  wire [2:0] _T_3174;
  reg [9:0] _T_3180;
  reg [31:0] _RAND_12;
  wire  _T_3182;
  wire  _T_3183;
  wire [1:0] _T_3184;
  wire [2:0] _T_3185;
  wire  _T_3187;
  wire  _T_3188;
  wire  _T_3190;
  reg [2:0] _T_3194;
  reg [31:0] _RAND_13;
  wire [2:0] _T_3195;
  wire [2:0] _T_3196;
  wire [5:0] _T_3197;
  wire [4:0] _T_3198;
  wire [5:0] _GEN_21;
  wire [5:0] _T_3199;
  wire [3:0] _T_3200;
  wire [5:0] _GEN_22;
  wire [5:0] _T_3201;
  wire [4:0] _T_3203;
  wire [5:0] _GEN_23;
  wire [5:0] _T_3204;
  wire [5:0] _GEN_24;
  wire [5:0] _T_3205;
  wire [2:0] _T_3206;
  wire [2:0] _T_3207;
  wire [2:0] _T_3208;
  wire [2:0] _T_3209;
  wire  _T_3211;
  wire  _T_3212;
  wire [2:0] _T_3213;
  wire [3:0] _GEN_25;
  wire [3:0] _T_3214;
  wire [2:0] _T_3215;
  wire [2:0] _T_3216;
  wire [4:0] _GEN_26;
  wire [4:0] _T_3217;
  wire [2:0] _T_3218;
  wire [2:0] _T_3219;
  wire [2:0] _GEN_3;
  wire  _T_3222;
  wire  _T_3223;
  wire  _T_3224;
  wire  _T_3233;
  wire  _T_3234;
  wire  _T_3235;
  wire  _T_3246;
  wire  _T_3247;
  wire  _T_3251;
  wire  _T_3256;
  wire  _T_3257;
  wire  _T_3259;
  wire  _T_3261;
  wire  _T_3262;
  wire  _T_3264;
  wire  _T_3265;
  wire  _T_3267;
  wire  _T_3268;
  wire  _T_3269;
  wire  _T_3271;
  wire  _T_3274;
  wire  _T_3275;
  wire  _T_3277;
  wire [9:0] _T_3279;
  wire [9:0] _T_3281;
  wire [9:0] _T_3283;
  wire [9:0] _T_3284;
  wire [9:0] _T_3285;
  wire  _T_3286;
  wire [9:0] _GEN_27;
  wire [10:0] _T_3287;
  wire [10:0] _T_3288;
  wire [9:0] _T_3289;
  wire [9:0] _T_3290;
  reg  _T_3312_0;
  reg [31:0] _RAND_14;
  reg  _T_3312_1;
  reg [31:0] _RAND_15;
  reg  _T_3312_2;
  reg [31:0] _RAND_16;
  wire  _T_3326_0;
  wire  _T_3326_1;
  wire  _T_3326_2;
  wire  _T_3336_0;
  wire  _T_3336_1;
  wire  _T_3336_2;
  wire  _T_3346;
  wire  _T_3347;
  wire  _T_3348;
  wire  _T_3353;
  wire  _T_3355;
  wire  _T_3357;
  wire  _T_3358;
  wire  _T_3359;
  wire  _T_3362;
  wire [32:0] _T_3364;
  wire [33:0] _T_3365;
  wire [8:0] _T_3366;
  wire [4:0] _T_3367;
  wire [13:0] _T_3368;
  wire [47:0] _T_3369;
  wire [47:0] _T_3371;
  wire [32:0] _T_3372;
  wire [33:0] _T_3373;
  wire [8:0] _T_3374;
  wire [4:0] _T_3375;
  wire [13:0] _T_3376;
  wire [47:0] _T_3377;
  wire [47:0] _T_3379;
  wire [32:0] _T_3380;
  wire [33:0] _T_3381;
  wire [8:0] _T_3382;
  wire [4:0] _T_3383;
  wire [13:0] _T_3384;
  wire [47:0] _T_3385;
  wire [47:0] _T_3387;
  wire [47:0] _T_3388;
  wire [47:0] _T_3389;
  wire  _T_3394;
  wire [31:0] _T_3395;
  wire [4:0] _T_3397;
  wire [3:0] _T_3398;
  wire [2:0] _T_3400;
  reg [9:0] _T_3404;
  reg [31:0] _RAND_17;
  wire  _T_3406;
  wire  _T_3407;
  wire [1:0] _T_3408;
  wire [2:0] _T_3409;
  wire  _T_3411;
  wire  _T_3412;
  wire  _T_3414;
  reg [2:0] _T_3418;
  reg [31:0] _RAND_18;
  wire [2:0] _T_3419;
  wire [2:0] _T_3420;
  wire [5:0] _T_3421;
  wire [4:0] _T_3422;
  wire [5:0] _GEN_28;
  wire [5:0] _T_3423;
  wire [3:0] _T_3424;
  wire [5:0] _GEN_29;
  wire [5:0] _T_3425;
  wire [4:0] _T_3427;
  wire [5:0] _GEN_30;
  wire [5:0] _T_3428;
  wire [5:0] _GEN_31;
  wire [5:0] _T_3429;
  wire [2:0] _T_3430;
  wire [2:0] _T_3431;
  wire [2:0] _T_3432;
  wire [2:0] _T_3433;
  wire  _T_3435;
  wire  _T_3436;
  wire [2:0] _T_3437;
  wire [3:0] _GEN_32;
  wire [3:0] _T_3438;
  wire [2:0] _T_3439;
  wire [2:0] _T_3440;
  wire [4:0] _GEN_33;
  wire [4:0] _T_3441;
  wire [2:0] _T_3442;
  wire [2:0] _T_3443;
  wire [2:0] _GEN_4;
  wire  _T_3446;
  wire  _T_3447;
  wire  _T_3448;
  wire  _T_3457;
  wire  _T_3458;
  wire  _T_3459;
  wire  _T_3470;
  wire  _T_3471;
  wire  _T_3475;
  wire  _T_3480;
  wire  _T_3481;
  wire  _T_3483;
  wire  _T_3485;
  wire  _T_3486;
  wire  _T_3488;
  wire  _T_3489;
  wire  _T_3491;
  wire  _T_3492;
  wire  _T_3493;
  wire  _T_3495;
  wire  _T_3498;
  wire  _T_3499;
  wire  _T_3501;
  wire [9:0] _T_3503;
  wire [9:0] _T_3505;
  wire [9:0] _T_3507;
  wire [9:0] _T_3508;
  wire [9:0] _T_3509;
  wire  _T_3510;
  wire [9:0] _GEN_34;
  wire [10:0] _T_3511;
  wire [10:0] _T_3512;
  wire [9:0] _T_3513;
  wire [9:0] _T_3514;
  reg  _T_3536_0;
  reg [31:0] _RAND_19;
  reg  _T_3536_1;
  reg [31:0] _RAND_20;
  reg  _T_3536_2;
  reg [31:0] _RAND_21;
  wire  _T_3550_0;
  wire  _T_3550_1;
  wire  _T_3550_2;
  wire  _T_3560_0;
  wire  _T_3560_1;
  wire  _T_3560_2;
  wire  _T_3570;
  wire  _T_3571;
  wire  _T_3572;
  wire  _T_3577;
  wire  _T_3579;
  wire  _T_3581;
  wire  _T_3582;
  wire  _T_3583;
  wire  _T_3586;
  wire [47:0] _T_3595;
  wire [47:0] _T_3603;
  wire [47:0] _T_3611;
  wire [47:0] _T_3612;
  wire [47:0] _T_3613;
  wire [4:0] _T_3621;
  wire [3:0] _T_3622;
  wire [2:0] _T_3624;
  assign io_in_1_a_ready = _T_2144;
  assign io_in_1_d_valid = _T_3586;
  assign io_in_1_d_bits_opcode = _T_3624;
  assign io_in_1_d_bits_size = _T_3622;
  assign io_in_1_d_bits_source = _T_504;
  assign io_in_0_a_ready = _T_2086;
  assign io_in_0_d_valid = _T_3362;
  assign io_in_0_d_bits_opcode = _T_3400;
  assign io_in_0_d_bits_size = _T_3398;
  assign io_in_0_d_bits_source = _T_495;
  assign io_in_0_d_bits_data = _T_3395;
  assign io_in_0_d_bits_error = _T_3394;
  assign io_out_2_a_valid = _T_3145;
  assign io_out_2_a_bits_opcode = _T_3174;
  assign io_out_2_a_bits_size = _T_3172;
  assign io_out_2_a_bits_source = _T_3171;
  assign io_out_2_d_ready = _T_2524;
  assign io_out_1_a_valid = _T_2967;
  assign io_out_1_a_bits_opcode = _T_2996;
  assign io_out_1_a_bits_size = _T_2994;
  assign io_out_1_a_bits_source = _T_2993;
  assign io_out_1_a_bits_address = _T_2992[30:0];
  assign io_out_1_a_bits_mask = _T_2991;
  assign io_out_1_a_bits_data = _T_2990;
  assign io_out_1_d_ready = _T_2480;
  assign io_out_0_a_valid = _T_2789;
  assign io_out_0_a_bits_opcode = _T_2818;
  assign io_out_0_a_bits_param = _T_2817;
  assign io_out_0_a_bits_size = _T_2816[2:0];
  assign io_out_0_a_bits_source = _T_2815;
  assign io_out_0_a_bits_address = _T_2814;
  assign io_out_0_a_bits_mask = _T_2813;
  assign io_out_0_a_bits_data = _T_2812;
  assign io_out_0_d_ready = _T_2436;
  assign in_1_a_bits_source = {{1'd0}, io_in_1_a_bits_source};
  assign _GEN_5 = {{4'd0}, io_in_0_a_bits_source};
  assign _T_494 = _GEN_5 | 5'h10;
  assign _T_495 = _T_3397[0];
  assign _T_504 = _T_3621[3:0];
  assign out_0_d_bits_size = {{1'd0}, io_out_0_d_bits_size};
  assign _T_908 = io_in_0_a_bits_address ^ 32'hc000000;
  assign _T_909 = {1'b0,$signed(_T_908)};
  assign _T_911 = $signed(_T_909) & $signed(33'shfc000000);
  assign _T_912 = $signed(_T_911);
  assign _T_914 = $signed(_T_912) == $signed(33'sh0);
  assign _T_916 = io_in_0_a_bits_address ^ 32'h2000000;
  assign _T_917 = {1'b0,$signed(_T_916)};
  assign _T_919 = $signed(_T_917) & $signed(33'shffff0000);
  assign _T_920 = $signed(_T_919);
  assign _T_922 = $signed(_T_920) == $signed(33'sh0);
  assign _T_925 = {1'b0,$signed(io_in_0_a_bits_address)};
  assign _T_927 = $signed(_T_925) & $signed(33'shffffd000);
  assign _T_928 = $signed(_T_927);
  assign _T_930 = $signed(_T_928) == $signed(33'sh0);
  assign _T_932 = io_in_0_a_bits_address ^ 32'h10000;
  assign _T_933 = {1'b0,$signed(_T_932)};
  assign _T_935 = $signed(_T_933) & $signed(33'shffff0000);
  assign _T_936 = $signed(_T_935);
  assign _T_938 = $signed(_T_936) == $signed(33'sh0);
  assign _T_940 = io_in_0_a_bits_address ^ 32'h80000000;
  assign _T_941 = {1'b0,$signed(_T_940)};
  assign _T_943 = $signed(_T_941) & $signed(33'shffffc000);
  assign _T_944 = $signed(_T_943);
  assign _T_946 = $signed(_T_944) == $signed(33'sh0);
  assign _T_947 = _T_914 | _T_922;
  assign _T_948 = _T_947 | _T_930;
  assign _T_949 = _T_948 | _T_938;
  assign _T_950 = _T_949 | _T_946;
  assign _T_952 = io_in_0_a_bits_address ^ 32'h60000000;
  assign _T_953 = {1'b0,$signed(_T_952)};
  assign _T_955 = $signed(_T_953) & $signed(33'she0000000);
  assign _T_956 = $signed(_T_955);
  assign _T_958 = $signed(_T_956) == $signed(33'sh0);
  assign _T_960 = io_in_0_a_bits_address ^ 32'h1000;
  assign _T_961 = {1'b0,$signed(_T_960)};
  assign _T_963 = $signed(_T_961) & $signed(33'shffffd000);
  assign _T_964 = $signed(_T_963);
  assign _T_966 = $signed(_T_964) == $signed(33'sh0);
  assign _T_976 = io_in_1_a_bits_address ^ 32'hc000000;
  assign _T_977 = {1'b0,$signed(_T_976)};
  assign _T_979 = $signed(_T_977) & $signed(33'shfc000000);
  assign _T_980 = $signed(_T_979);
  assign _T_982 = $signed(_T_980) == $signed(33'sh0);
  assign _T_984 = io_in_1_a_bits_address ^ 32'h2000000;
  assign _T_985 = {1'b0,$signed(_T_984)};
  assign _T_987 = $signed(_T_985) & $signed(33'shffff0000);
  assign _T_988 = $signed(_T_987);
  assign _T_990 = $signed(_T_988) == $signed(33'sh0);
  assign _T_993 = {1'b0,$signed(io_in_1_a_bits_address)};
  assign _T_995 = $signed(_T_993) & $signed(33'shffffd000);
  assign _T_996 = $signed(_T_995);
  assign _T_998 = $signed(_T_996) == $signed(33'sh0);
  assign _T_1000 = io_in_1_a_bits_address ^ 32'h10000;
  assign _T_1001 = {1'b0,$signed(_T_1000)};
  assign _T_1003 = $signed(_T_1001) & $signed(33'shffff0000);
  assign _T_1004 = $signed(_T_1003);
  assign _T_1006 = $signed(_T_1004) == $signed(33'sh0);
  assign _T_1008 = io_in_1_a_bits_address ^ 32'h80000000;
  assign _T_1009 = {1'b0,$signed(_T_1008)};
  assign _T_1011 = $signed(_T_1009) & $signed(33'shffffc000);
  assign _T_1012 = $signed(_T_1011);
  assign _T_1014 = $signed(_T_1012) == $signed(33'sh0);
  assign _T_1015 = _T_982 | _T_990;
  assign _T_1016 = _T_1015 | _T_998;
  assign _T_1017 = _T_1016 | _T_1006;
  assign _T_1018 = _T_1017 | _T_1014;
  assign _T_1020 = io_in_1_a_bits_address ^ 32'h60000000;
  assign _T_1021 = {1'b0,$signed(_T_1020)};
  assign _T_1023 = $signed(_T_1021) & $signed(33'she0000000);
  assign _T_1024 = $signed(_T_1023);
  assign _T_1026 = $signed(_T_1024) == $signed(33'sh0);
  assign _T_1028 = io_in_1_a_bits_address ^ 32'h1000;
  assign _T_1029 = {1'b0,$signed(_T_1028)};
  assign _T_1031 = $signed(_T_1029) & $signed(33'shffffd000);
  assign _T_1032 = $signed(_T_1031);
  assign _T_1034 = $signed(_T_1032) == $signed(33'sh0);
  assign _T_1576 = io_out_0_d_bits_source[4:1];
  assign _T_1578 = _T_1576 == 4'h8;
  assign _T_1588 = io_out_0_d_bits_source[4:4];
  assign _T_1590 = _T_1588 == 1'h0;
  assign _T_1607 = io_out_1_d_bits_source[4:1];
  assign _T_1609 = _T_1607 == 4'h8;
  assign _T_1619 = io_out_1_d_bits_source[4:4];
  assign _T_1621 = _T_1619 == 1'h0;
  assign _T_1638 = io_out_2_d_bits_source[4:1];
  assign _T_1640 = _T_1638 == 4'h8;
  assign _T_1650 = io_out_2_d_bits_source[4:4];
  assign _T_1652 = _T_1650 == 1'h0;
  assign _T_1894 = 27'hfff << io_in_0_a_bits_size;
  assign _T_1895 = _T_1894[11:0];
  assign _T_1896 = ~ _T_1895;
  assign _T_1897 = _T_1896[11:2];
  assign _T_1898 = io_in_0_a_bits_opcode[2];
  assign _T_1900 = _T_1898 == 1'h0;
  assign _T_1902 = _T_1900 ? _T_1897 : 10'h0;
  assign _T_1905 = 27'hfff << io_in_1_a_bits_size;
  assign _T_1906 = _T_1905[11:0];
  assign _T_1907 = ~ _T_1906;
  assign _T_1908 = _T_1907[11:2];
  assign _T_1909 = io_in_1_a_bits_opcode[2];
  assign _T_1911 = _T_1909 == 1'h0;
  assign _T_1913 = _T_1911 ? _T_1908 : 10'h0;
  assign _T_1991 = 21'h3f << out_0_d_bits_size;
  assign _T_1992 = _T_1991[5:0];
  assign _T_1993 = ~ _T_1992;
  assign _T_1994 = _T_1993[5:2];
  assign _T_1995 = io_out_0_d_bits_opcode[0];
  assign _T_1997 = _T_1995 ? _T_1994 : 4'h0;
  assign _T_2000 = 23'hff << io_out_1_d_bits_size;
  assign _T_2001 = _T_2000[7:0];
  assign _T_2002 = ~ _T_2001;
  assign _T_2003 = _T_2002[7:2];
  assign _T_2004 = io_out_1_d_bits_opcode[0];
  assign _T_2006 = _T_2004 ? _T_2003 : 6'h0;
  assign _T_2009 = 27'hfff << io_out_2_d_bits_size;
  assign _T_2010 = _T_2009[11:0];
  assign _T_2011 = ~ _T_2010;
  assign _T_2012 = _T_2011[11:2];
  assign _T_2013 = io_out_2_d_bits_opcode[0];
  assign _T_2015 = _T_2013 ? _T_2012 : 10'h0;
  assign beatsDO_0 = {{6'd0}, _T_1997};
  assign beatsDO_1 = {{4'd0}, _T_2006};
  assign _T_2075 = io_in_0_a_valid & _T_950;
  assign _T_2076 = io_in_0_a_valid & _T_958;
  assign _T_2077 = io_in_0_a_valid & _T_966;
  assign _T_2080 = _T_950 ? _T_2778 : 1'h0;
  assign _T_2082 = _T_958 ? _T_2956 : 1'h0;
  assign _T_2084 = _T_966 ? _T_3134 : 1'h0;
  assign _T_2085 = _T_2080 | _T_2082;
  assign _T_2086 = _T_2085 | _T_2084;
  assign _T_2133 = io_in_1_a_valid & _T_1018;
  assign _T_2134 = io_in_1_a_valid & _T_1026;
  assign _T_2135 = io_in_1_a_valid & _T_1034;
  assign _T_2138 = _T_1018 ? _T_2779 : 1'h0;
  assign _T_2140 = _T_1026 ? _T_2957 : 1'h0;
  assign _T_2142 = _T_1034 ? _T_3135 : 1'h0;
  assign _T_2143 = _T_2138 | _T_2140;
  assign _T_2144 = _T_2143 | _T_2142;
  assign _T_2429 = io_out_0_d_valid & _T_1578;
  assign _T_2430 = io_out_0_d_valid & _T_1590;
  assign _T_2433 = _T_1578 ? _T_3346 : 1'h0;
  assign _T_2435 = _T_1590 ? _T_3570 : 1'h0;
  assign _T_2436 = _T_2433 | _T_2435;
  assign _T_2473 = io_out_1_d_valid & _T_1609;
  assign _T_2474 = io_out_1_d_valid & _T_1621;
  assign _T_2477 = _T_1609 ? _T_3347 : 1'h0;
  assign _T_2479 = _T_1621 ? _T_3571 : 1'h0;
  assign _T_2480 = _T_2477 | _T_2479;
  assign _T_2517 = io_out_2_d_valid & _T_1640;
  assign _T_2518 = io_out_2_d_valid & _T_1652;
  assign _T_2521 = _T_1640 ? _T_3348 : 1'h0;
  assign _T_2523 = _T_1652 ? _T_3572 : 1'h0;
  assign _T_2524 = _T_2521 | _T_2523;
  assign _T_2647 = _T_2645 == 10'h0;
  assign _T_2648 = _T_2647 & io_out_0_a_ready;
  assign _T_2649 = {_T_2133,_T_2075};
  assign _T_2651 = _T_2649 == _T_2649;
  assign _T_2652 = _T_2651 | reset;
  assign _T_2654 = _T_2652 == 1'h0;
  assign _T_2659 = ~ _T_2658;
  assign _T_2660 = _T_2649 & _T_2659;
  assign _T_2661 = {_T_2660,_T_2649};
  assign _T_2662 = _T_2661[3:1];
  assign _GEN_6 = {{1'd0}, _T_2662};
  assign _T_2663 = _T_2661 | _GEN_6;
  assign _T_2665 = _T_2663[3:1];
  assign _GEN_7 = {{2'd0}, _T_2658};
  assign _T_2666 = _GEN_7 << 2;
  assign _GEN_8 = {{1'd0}, _T_2665};
  assign _T_2667 = _GEN_8 | _T_2666;
  assign _T_2668 = _T_2667[3:2];
  assign _T_2669 = _T_2667[1:0];
  assign _T_2670 = _T_2668 & _T_2669;
  assign _T_2671 = ~ _T_2670;
  assign _T_2673 = _T_2649 != 2'h0;
  assign _T_2674 = _T_2648 & _T_2673;
  assign _T_2675 = _T_2671 & _T_2649;
  assign _GEN_9 = {{1'd0}, _T_2675};
  assign _T_2676 = _GEN_9 << 1;
  assign _T_2677 = _T_2676[1:0];
  assign _T_2678 = _T_2675 | _T_2677;
  assign _GEN_0 = _T_2674 ? _T_2678 : _T_2658;
  assign _T_2681 = _T_2671[0];
  assign _T_2682 = _T_2671[1];
  assign _T_2690 = _T_2681 & _T_2075;
  assign _T_2691 = _T_2682 & _T_2133;
  assign _T_2701 = _T_2690 | _T_2691;
  assign _T_2705 = _T_2690 == 1'h0;
  assign _T_2710 = _T_2691 == 1'h0;
  assign _T_2711 = _T_2705 | _T_2710;
  assign _T_2713 = _T_2711 | reset;
  assign _T_2715 = _T_2713 == 1'h0;
  assign _T_2716 = _T_2075 | _T_2133;
  assign _T_2718 = _T_2716 == 1'h0;
  assign _T_2720 = _T_2718 | _T_2701;
  assign _T_2721 = _T_2720 | reset;
  assign _T_2723 = _T_2721 == 1'h0;
  assign _T_2725 = _T_2690 ? _T_1902 : 10'h0;
  assign _T_2727 = _T_2691 ? _T_1913 : 10'h0;
  assign _T_2728 = _T_2725 | _T_2727;
  assign _T_2729 = io_out_0_a_ready & _T_2789;
  assign _GEN_10 = {{9'd0}, _T_2729};
  assign _T_2730 = _T_2645 - _GEN_10;
  assign _T_2731 = $unsigned(_T_2730);
  assign _T_2732 = _T_2731[9:0];
  assign _T_2733 = _T_2648 ? _T_2728 : _T_2732;
  assign _T_2762_0 = _T_2647 ? _T_2690 : _T_2751_0;
  assign _T_2762_1 = _T_2647 ? _T_2691 : _T_2751_1;
  assign _T_2770_0 = _T_2647 ? _T_2681 : _T_2751_0;
  assign _T_2770_1 = _T_2647 ? _T_2682 : _T_2751_1;
  assign _T_2778 = io_out_0_a_ready & _T_2770_0;
  assign _T_2779 = io_out_0_a_ready & _T_2770_1;
  assign _T_2783 = _T_2751_0 ? _T_2075 : 1'h0;
  assign _T_2785 = _T_2751_1 ? _T_2133 : 1'h0;
  assign _T_2786 = _T_2783 | _T_2785;
  assign _T_2789 = _T_2647 ? _T_2716 : _T_2786;
  assign _T_2791 = {io_in_0_a_bits_address,io_in_0_a_bits_mask};
  assign _T_2792 = {_T_2791,io_in_0_a_bits_data};
  assign _T_2793 = {io_in_0_a_bits_size,_T_494};
  assign _T_2794 = {io_in_0_a_bits_opcode,io_in_0_a_bits_param};
  assign _T_2795 = {_T_2794,_T_2793};
  assign _T_2796 = {_T_2795,_T_2792};
  assign _T_2798 = _T_2762_0 ? _T_2796 : 83'h0;
  assign _T_2799 = {io_in_1_a_bits_address,io_in_1_a_bits_mask};
  assign _T_2800 = {_T_2799,io_in_1_a_bits_data};
  assign _T_2801 = {io_in_1_a_bits_size,in_1_a_bits_source};
  assign _T_2802 = {io_in_1_a_bits_opcode,io_in_1_a_bits_param};
  assign _T_2803 = {_T_2802,_T_2801};
  assign _T_2804 = {_T_2803,_T_2800};
  assign _T_2806 = _T_2762_1 ? _T_2804 : 83'h0;
  assign _T_2807 = _T_2798 | _T_2806;
  assign _T_2812 = _T_2807[31:0];
  assign _T_2813 = _T_2807[35:32];
  assign _T_2814 = _T_2807[67:36];
  assign _T_2815 = _T_2807[72:68];
  assign _T_2816 = _T_2807[76:73];
  assign _T_2817 = _T_2807[79:77];
  assign _T_2818 = _T_2807[82:80];
  assign _T_2825 = _T_2823 == 10'h0;
  assign _T_2826 = _T_2825 & io_out_1_a_ready;
  assign _T_2827 = {_T_2134,_T_2076};
  assign _T_2829 = _T_2827 == _T_2827;
  assign _T_2830 = _T_2829 | reset;
  assign _T_2832 = _T_2830 == 1'h0;
  assign _T_2837 = ~ _T_2836;
  assign _T_2838 = _T_2827 & _T_2837;
  assign _T_2839 = {_T_2838,_T_2827};
  assign _T_2840 = _T_2839[3:1];
  assign _GEN_11 = {{1'd0}, _T_2840};
  assign _T_2841 = _T_2839 | _GEN_11;
  assign _T_2843 = _T_2841[3:1];
  assign _GEN_12 = {{2'd0}, _T_2836};
  assign _T_2844 = _GEN_12 << 2;
  assign _GEN_13 = {{1'd0}, _T_2843};
  assign _T_2845 = _GEN_13 | _T_2844;
  assign _T_2846 = _T_2845[3:2];
  assign _T_2847 = _T_2845[1:0];
  assign _T_2848 = _T_2846 & _T_2847;
  assign _T_2849 = ~ _T_2848;
  assign _T_2851 = _T_2827 != 2'h0;
  assign _T_2852 = _T_2826 & _T_2851;
  assign _T_2853 = _T_2849 & _T_2827;
  assign _GEN_14 = {{1'd0}, _T_2853};
  assign _T_2854 = _GEN_14 << 1;
  assign _T_2855 = _T_2854[1:0];
  assign _T_2856 = _T_2853 | _T_2855;
  assign _GEN_1 = _T_2852 ? _T_2856 : _T_2836;
  assign _T_2859 = _T_2849[0];
  assign _T_2860 = _T_2849[1];
  assign _T_2868 = _T_2859 & _T_2076;
  assign _T_2869 = _T_2860 & _T_2134;
  assign _T_2879 = _T_2868 | _T_2869;
  assign _T_2883 = _T_2868 == 1'h0;
  assign _T_2888 = _T_2869 == 1'h0;
  assign _T_2889 = _T_2883 | _T_2888;
  assign _T_2891 = _T_2889 | reset;
  assign _T_2893 = _T_2891 == 1'h0;
  assign _T_2894 = _T_2076 | _T_2134;
  assign _T_2896 = _T_2894 == 1'h0;
  assign _T_2898 = _T_2896 | _T_2879;
  assign _T_2899 = _T_2898 | reset;
  assign _T_2901 = _T_2899 == 1'h0;
  assign _T_2903 = _T_2868 ? _T_1902 : 10'h0;
  assign _T_2905 = _T_2869 ? _T_1913 : 10'h0;
  assign _T_2906 = _T_2903 | _T_2905;
  assign _T_2907 = io_out_1_a_ready & _T_2967;
  assign _GEN_15 = {{9'd0}, _T_2907};
  assign _T_2908 = _T_2823 - _GEN_15;
  assign _T_2909 = $unsigned(_T_2908);
  assign _T_2910 = _T_2909[9:0];
  assign _T_2911 = _T_2826 ? _T_2906 : _T_2910;
  assign _T_2940_0 = _T_2825 ? _T_2868 : _T_2929_0;
  assign _T_2940_1 = _T_2825 ? _T_2869 : _T_2929_1;
  assign _T_2948_0 = _T_2825 ? _T_2859 : _T_2929_0;
  assign _T_2948_1 = _T_2825 ? _T_2860 : _T_2929_1;
  assign _T_2956 = io_out_1_a_ready & _T_2948_0;
  assign _T_2957 = io_out_1_a_ready & _T_2948_1;
  assign _T_2961 = _T_2929_0 ? _T_2076 : 1'h0;
  assign _T_2963 = _T_2929_1 ? _T_2134 : 1'h0;
  assign _T_2964 = _T_2961 | _T_2963;
  assign _T_2967 = _T_2825 ? _T_2894 : _T_2964;
  assign _T_2976 = _T_2940_0 ? _T_2796 : 83'h0;
  assign _T_2984 = _T_2940_1 ? _T_2804 : 83'h0;
  assign _T_2985 = _T_2976 | _T_2984;
  assign _T_2990 = _T_2985[31:0];
  assign _T_2991 = _T_2985[35:32];
  assign _T_2992 = _T_2985[67:36];
  assign _T_2993 = _T_2985[72:68];
  assign _T_2994 = _T_2985[76:73];
  assign _T_2996 = _T_2985[82:80];
  assign _T_3003 = _T_3001 == 10'h0;
  assign _T_3004 = _T_3003 & io_out_2_a_ready;
  assign _T_3005 = {_T_2135,_T_2077};
  assign _T_3007 = _T_3005 == _T_3005;
  assign _T_3008 = _T_3007 | reset;
  assign _T_3010 = _T_3008 == 1'h0;
  assign _T_3015 = ~ _T_3014;
  assign _T_3016 = _T_3005 & _T_3015;
  assign _T_3017 = {_T_3016,_T_3005};
  assign _T_3018 = _T_3017[3:1];
  assign _GEN_16 = {{1'd0}, _T_3018};
  assign _T_3019 = _T_3017 | _GEN_16;
  assign _T_3021 = _T_3019[3:1];
  assign _GEN_17 = {{2'd0}, _T_3014};
  assign _T_3022 = _GEN_17 << 2;
  assign _GEN_18 = {{1'd0}, _T_3021};
  assign _T_3023 = _GEN_18 | _T_3022;
  assign _T_3024 = _T_3023[3:2];
  assign _T_3025 = _T_3023[1:0];
  assign _T_3026 = _T_3024 & _T_3025;
  assign _T_3027 = ~ _T_3026;
  assign _T_3029 = _T_3005 != 2'h0;
  assign _T_3030 = _T_3004 & _T_3029;
  assign _T_3031 = _T_3027 & _T_3005;
  assign _GEN_19 = {{1'd0}, _T_3031};
  assign _T_3032 = _GEN_19 << 1;
  assign _T_3033 = _T_3032[1:0];
  assign _T_3034 = _T_3031 | _T_3033;
  assign _GEN_2 = _T_3030 ? _T_3034 : _T_3014;
  assign _T_3037 = _T_3027[0];
  assign _T_3038 = _T_3027[1];
  assign _T_3046 = _T_3037 & _T_2077;
  assign _T_3047 = _T_3038 & _T_2135;
  assign _T_3057 = _T_3046 | _T_3047;
  assign _T_3061 = _T_3046 == 1'h0;
  assign _T_3066 = _T_3047 == 1'h0;
  assign _T_3067 = _T_3061 | _T_3066;
  assign _T_3069 = _T_3067 | reset;
  assign _T_3071 = _T_3069 == 1'h0;
  assign _T_3072 = _T_2077 | _T_2135;
  assign _T_3074 = _T_3072 == 1'h0;
  assign _T_3076 = _T_3074 | _T_3057;
  assign _T_3077 = _T_3076 | reset;
  assign _T_3079 = _T_3077 == 1'h0;
  assign _T_3081 = _T_3046 ? _T_1902 : 10'h0;
  assign _T_3083 = _T_3047 ? _T_1913 : 10'h0;
  assign _T_3084 = _T_3081 | _T_3083;
  assign _T_3085 = io_out_2_a_ready & _T_3145;
  assign _GEN_20 = {{9'd0}, _T_3085};
  assign _T_3086 = _T_3001 - _GEN_20;
  assign _T_3087 = $unsigned(_T_3086);
  assign _T_3088 = _T_3087[9:0];
  assign _T_3089 = _T_3004 ? _T_3084 : _T_3088;
  assign _T_3118_0 = _T_3003 ? _T_3046 : _T_3107_0;
  assign _T_3118_1 = _T_3003 ? _T_3047 : _T_3107_1;
  assign _T_3126_0 = _T_3003 ? _T_3037 : _T_3107_0;
  assign _T_3126_1 = _T_3003 ? _T_3038 : _T_3107_1;
  assign _T_3134 = io_out_2_a_ready & _T_3126_0;
  assign _T_3135 = io_out_2_a_ready & _T_3126_1;
  assign _T_3139 = _T_3107_0 ? _T_2077 : 1'h0;
  assign _T_3141 = _T_3107_1 ? _T_2135 : 1'h0;
  assign _T_3142 = _T_3139 | _T_3141;
  assign _T_3145 = _T_3003 ? _T_3072 : _T_3142;
  assign _T_3154 = _T_3118_0 ? _T_2796 : 83'h0;
  assign _T_3162 = _T_3118_1 ? _T_2804 : 83'h0;
  assign _T_3163 = _T_3154 | _T_3162;
  assign _T_3171 = _T_3163[72:68];
  assign _T_3172 = _T_3163[76:73];
  assign _T_3174 = _T_3163[82:80];
  assign _T_3182 = _T_3180 == 10'h0;
  assign _T_3183 = _T_3182 & io_in_0_d_ready;
  assign _T_3184 = {_T_2517,_T_2473};
  assign _T_3185 = {_T_3184,_T_2429};
  assign _T_3187 = _T_3185 == _T_3185;
  assign _T_3188 = _T_3187 | reset;
  assign _T_3190 = _T_3188 == 1'h0;
  assign _T_3195 = ~ _T_3194;
  assign _T_3196 = _T_3185 & _T_3195;
  assign _T_3197 = {_T_3196,_T_3185};
  assign _T_3198 = _T_3197[5:1];
  assign _GEN_21 = {{1'd0}, _T_3198};
  assign _T_3199 = _T_3197 | _GEN_21;
  assign _T_3200 = _T_3199[5:2];
  assign _GEN_22 = {{2'd0}, _T_3200};
  assign _T_3201 = _T_3199 | _GEN_22;
  assign _T_3203 = _T_3201[5:1];
  assign _GEN_23 = {{3'd0}, _T_3194};
  assign _T_3204 = _GEN_23 << 3;
  assign _GEN_24 = {{1'd0}, _T_3203};
  assign _T_3205 = _GEN_24 | _T_3204;
  assign _T_3206 = _T_3205[5:3];
  assign _T_3207 = _T_3205[2:0];
  assign _T_3208 = _T_3206 & _T_3207;
  assign _T_3209 = ~ _T_3208;
  assign _T_3211 = _T_3185 != 3'h0;
  assign _T_3212 = _T_3183 & _T_3211;
  assign _T_3213 = _T_3209 & _T_3185;
  assign _GEN_25 = {{1'd0}, _T_3213};
  assign _T_3214 = _GEN_25 << 1;
  assign _T_3215 = _T_3214[2:0];
  assign _T_3216 = _T_3213 | _T_3215;
  assign _GEN_26 = {{2'd0}, _T_3216};
  assign _T_3217 = _GEN_26 << 2;
  assign _T_3218 = _T_3217[2:0];
  assign _T_3219 = _T_3216 | _T_3218;
  assign _GEN_3 = _T_3212 ? _T_3219 : _T_3194;
  assign _T_3222 = _T_3209[0];
  assign _T_3223 = _T_3209[1];
  assign _T_3224 = _T_3209[2];
  assign _T_3233 = _T_3222 & _T_2429;
  assign _T_3234 = _T_3223 & _T_2473;
  assign _T_3235 = _T_3224 & _T_2517;
  assign _T_3246 = _T_3233 | _T_3234;
  assign _T_3247 = _T_3246 | _T_3235;
  assign _T_3251 = _T_3233 == 1'h0;
  assign _T_3256 = _T_3234 == 1'h0;
  assign _T_3257 = _T_3251 | _T_3256;
  assign _T_3259 = _T_3246 == 1'h0;
  assign _T_3261 = _T_3235 == 1'h0;
  assign _T_3262 = _T_3259 | _T_3261;
  assign _T_3264 = _T_3257 & _T_3262;
  assign _T_3265 = _T_3264 | reset;
  assign _T_3267 = _T_3265 == 1'h0;
  assign _T_3268 = _T_2429 | _T_2473;
  assign _T_3269 = _T_3268 | _T_2517;
  assign _T_3271 = _T_3269 == 1'h0;
  assign _T_3274 = _T_3271 | _T_3247;
  assign _T_3275 = _T_3274 | reset;
  assign _T_3277 = _T_3275 == 1'h0;
  assign _T_3279 = _T_3233 ? beatsDO_0 : 10'h0;
  assign _T_3281 = _T_3234 ? beatsDO_1 : 10'h0;
  assign _T_3283 = _T_3235 ? _T_2015 : 10'h0;
  assign _T_3284 = _T_3279 | _T_3281;
  assign _T_3285 = _T_3284 | _T_3283;
  assign _T_3286 = io_in_0_d_ready & _T_3362;
  assign _GEN_27 = {{9'd0}, _T_3286};
  assign _T_3287 = _T_3180 - _GEN_27;
  assign _T_3288 = $unsigned(_T_3287);
  assign _T_3289 = _T_3288[9:0];
  assign _T_3290 = _T_3183 ? _T_3285 : _T_3289;
  assign _T_3326_0 = _T_3182 ? _T_3233 : _T_3312_0;
  assign _T_3326_1 = _T_3182 ? _T_3234 : _T_3312_1;
  assign _T_3326_2 = _T_3182 ? _T_3235 : _T_3312_2;
  assign _T_3336_0 = _T_3182 ? _T_3222 : _T_3312_0;
  assign _T_3336_1 = _T_3182 ? _T_3223 : _T_3312_1;
  assign _T_3336_2 = _T_3182 ? _T_3224 : _T_3312_2;
  assign _T_3346 = io_in_0_d_ready & _T_3336_0;
  assign _T_3347 = io_in_0_d_ready & _T_3336_1;
  assign _T_3348 = io_in_0_d_ready & _T_3336_2;
  assign _T_3353 = _T_3312_0 ? _T_2429 : 1'h0;
  assign _T_3355 = _T_3312_1 ? _T_2473 : 1'h0;
  assign _T_3357 = _T_3312_2 ? _T_2517 : 1'h0;
  assign _T_3358 = _T_3353 | _T_3355;
  assign _T_3359 = _T_3358 | _T_3357;
  assign _T_3362 = _T_3182 ? _T_3269 : _T_3359;
  assign _T_3364 = {io_out_0_d_bits_sink,io_out_0_d_bits_data};
  assign _T_3365 = {_T_3364,io_out_0_d_bits_error};
  assign _T_3366 = {out_0_d_bits_size,io_out_0_d_bits_source};
  assign _T_3367 = {io_out_0_d_bits_opcode,io_out_0_d_bits_param};
  assign _T_3368 = {_T_3367,_T_3366};
  assign _T_3369 = {_T_3368,_T_3365};
  assign _T_3371 = _T_3326_0 ? _T_3369 : 48'h0;
  assign _T_3372 = {io_out_1_d_bits_sink,io_out_1_d_bits_data};
  assign _T_3373 = {_T_3372,io_out_1_d_bits_error};
  assign _T_3374 = {io_out_1_d_bits_size,io_out_1_d_bits_source};
  assign _T_3375 = {io_out_1_d_bits_opcode,io_out_1_d_bits_param};
  assign _T_3376 = {_T_3375,_T_3374};
  assign _T_3377 = {_T_3376,_T_3373};
  assign _T_3379 = _T_3326_1 ? _T_3377 : 48'h0;
  assign _T_3380 = {io_out_2_d_bits_sink,io_out_2_d_bits_data};
  assign _T_3381 = {_T_3380,io_out_2_d_bits_error};
  assign _T_3382 = {io_out_2_d_bits_size,io_out_2_d_bits_source};
  assign _T_3383 = {io_out_2_d_bits_opcode,io_out_2_d_bits_param};
  assign _T_3384 = {_T_3383,_T_3382};
  assign _T_3385 = {_T_3384,_T_3381};
  assign _T_3387 = _T_3326_2 ? _T_3385 : 48'h0;
  assign _T_3388 = _T_3371 | _T_3379;
  assign _T_3389 = _T_3388 | _T_3387;
  assign _T_3394 = _T_3389[0];
  assign _T_3395 = _T_3389[32:1];
  assign _T_3397 = _T_3389[38:34];
  assign _T_3398 = _T_3389[42:39];
  assign _T_3400 = _T_3389[47:45];
  assign _T_3406 = _T_3404 == 10'h0;
  assign _T_3407 = _T_3406 & io_in_1_d_ready;
  assign _T_3408 = {_T_2518,_T_2474};
  assign _T_3409 = {_T_3408,_T_2430};
  assign _T_3411 = _T_3409 == _T_3409;
  assign _T_3412 = _T_3411 | reset;
  assign _T_3414 = _T_3412 == 1'h0;
  assign _T_3419 = ~ _T_3418;
  assign _T_3420 = _T_3409 & _T_3419;
  assign _T_3421 = {_T_3420,_T_3409};
  assign _T_3422 = _T_3421[5:1];
  assign _GEN_28 = {{1'd0}, _T_3422};
  assign _T_3423 = _T_3421 | _GEN_28;
  assign _T_3424 = _T_3423[5:2];
  assign _GEN_29 = {{2'd0}, _T_3424};
  assign _T_3425 = _T_3423 | _GEN_29;
  assign _T_3427 = _T_3425[5:1];
  assign _GEN_30 = {{3'd0}, _T_3418};
  assign _T_3428 = _GEN_30 << 3;
  assign _GEN_31 = {{1'd0}, _T_3427};
  assign _T_3429 = _GEN_31 | _T_3428;
  assign _T_3430 = _T_3429[5:3];
  assign _T_3431 = _T_3429[2:0];
  assign _T_3432 = _T_3430 & _T_3431;
  assign _T_3433 = ~ _T_3432;
  assign _T_3435 = _T_3409 != 3'h0;
  assign _T_3436 = _T_3407 & _T_3435;
  assign _T_3437 = _T_3433 & _T_3409;
  assign _GEN_32 = {{1'd0}, _T_3437};
  assign _T_3438 = _GEN_32 << 1;
  assign _T_3439 = _T_3438[2:0];
  assign _T_3440 = _T_3437 | _T_3439;
  assign _GEN_33 = {{2'd0}, _T_3440};
  assign _T_3441 = _GEN_33 << 2;
  assign _T_3442 = _T_3441[2:0];
  assign _T_3443 = _T_3440 | _T_3442;
  assign _GEN_4 = _T_3436 ? _T_3443 : _T_3418;
  assign _T_3446 = _T_3433[0];
  assign _T_3447 = _T_3433[1];
  assign _T_3448 = _T_3433[2];
  assign _T_3457 = _T_3446 & _T_2430;
  assign _T_3458 = _T_3447 & _T_2474;
  assign _T_3459 = _T_3448 & _T_2518;
  assign _T_3470 = _T_3457 | _T_3458;
  assign _T_3471 = _T_3470 | _T_3459;
  assign _T_3475 = _T_3457 == 1'h0;
  assign _T_3480 = _T_3458 == 1'h0;
  assign _T_3481 = _T_3475 | _T_3480;
  assign _T_3483 = _T_3470 == 1'h0;
  assign _T_3485 = _T_3459 == 1'h0;
  assign _T_3486 = _T_3483 | _T_3485;
  assign _T_3488 = _T_3481 & _T_3486;
  assign _T_3489 = _T_3488 | reset;
  assign _T_3491 = _T_3489 == 1'h0;
  assign _T_3492 = _T_2430 | _T_2474;
  assign _T_3493 = _T_3492 | _T_2518;
  assign _T_3495 = _T_3493 == 1'h0;
  assign _T_3498 = _T_3495 | _T_3471;
  assign _T_3499 = _T_3498 | reset;
  assign _T_3501 = _T_3499 == 1'h0;
  assign _T_3503 = _T_3457 ? beatsDO_0 : 10'h0;
  assign _T_3505 = _T_3458 ? beatsDO_1 : 10'h0;
  assign _T_3507 = _T_3459 ? _T_2015 : 10'h0;
  assign _T_3508 = _T_3503 | _T_3505;
  assign _T_3509 = _T_3508 | _T_3507;
  assign _T_3510 = io_in_1_d_ready & _T_3586;
  assign _GEN_34 = {{9'd0}, _T_3510};
  assign _T_3511 = _T_3404 - _GEN_34;
  assign _T_3512 = $unsigned(_T_3511);
  assign _T_3513 = _T_3512[9:0];
  assign _T_3514 = _T_3407 ? _T_3509 : _T_3513;
  assign _T_3550_0 = _T_3406 ? _T_3457 : _T_3536_0;
  assign _T_3550_1 = _T_3406 ? _T_3458 : _T_3536_1;
  assign _T_3550_2 = _T_3406 ? _T_3459 : _T_3536_2;
  assign _T_3560_0 = _T_3406 ? _T_3446 : _T_3536_0;
  assign _T_3560_1 = _T_3406 ? _T_3447 : _T_3536_1;
  assign _T_3560_2 = _T_3406 ? _T_3448 : _T_3536_2;
  assign _T_3570 = io_in_1_d_ready & _T_3560_0;
  assign _T_3571 = io_in_1_d_ready & _T_3560_1;
  assign _T_3572 = io_in_1_d_ready & _T_3560_2;
  assign _T_3577 = _T_3536_0 ? _T_2430 : 1'h0;
  assign _T_3579 = _T_3536_1 ? _T_2474 : 1'h0;
  assign _T_3581 = _T_3536_2 ? _T_2518 : 1'h0;
  assign _T_3582 = _T_3577 | _T_3579;
  assign _T_3583 = _T_3582 | _T_3581;
  assign _T_3586 = _T_3406 ? _T_3493 : _T_3583;
  assign _T_3595 = _T_3550_0 ? _T_3369 : 48'h0;
  assign _T_3603 = _T_3550_1 ? _T_3377 : 48'h0;
  assign _T_3611 = _T_3550_2 ? _T_3385 : 48'h0;
  assign _T_3612 = _T_3595 | _T_3603;
  assign _T_3613 = _T_3612 | _T_3611;
  assign _T_3621 = _T_3613[38:34];
  assign _T_3622 = _T_3613[42:39];
  assign _T_3624 = _T_3613[47:45];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_2645 = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_2658 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_2751_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_2751_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_2823 = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_2836 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_2929_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_2929_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_3001 = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_3014 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_3107_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_3107_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_3180 = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_3194 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_3312_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_3312_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_3312_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_3404 = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_3418 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_3536_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_3536_1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_3536_2 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_2645 <= 10'h0;
    end else begin
      if (_T_2648) begin
        _T_2645 <= _T_2728;
      end else begin
        _T_2645 <= _T_2732;
      end
    end
    if (reset) begin
      _T_2658 <= 2'h3;
    end else begin
      if (_T_2674) begin
        _T_2658 <= _T_2678;
      end
    end
    if (reset) begin
      _T_2751_0 <= 1'h0;
    end else begin
      if (_T_2647) begin
        _T_2751_0 <= _T_2690;
      end
    end
    if (reset) begin
      _T_2751_1 <= 1'h0;
    end else begin
      if (_T_2647) begin
        _T_2751_1 <= _T_2691;
      end
    end
    if (reset) begin
      _T_2823 <= 10'h0;
    end else begin
      if (_T_2826) begin
        _T_2823 <= _T_2906;
      end else begin
        _T_2823 <= _T_2910;
      end
    end
    if (reset) begin
      _T_2836 <= 2'h3;
    end else begin
      if (_T_2852) begin
        _T_2836 <= _T_2856;
      end
    end
    if (reset) begin
      _T_2929_0 <= 1'h0;
    end else begin
      if (_T_2825) begin
        _T_2929_0 <= _T_2868;
      end
    end
    if (reset) begin
      _T_2929_1 <= 1'h0;
    end else begin
      if (_T_2825) begin
        _T_2929_1 <= _T_2869;
      end
    end
    if (reset) begin
      _T_3001 <= 10'h0;
    end else begin
      if (_T_3004) begin
        _T_3001 <= _T_3084;
      end else begin
        _T_3001 <= _T_3088;
      end
    end
    if (reset) begin
      _T_3014 <= 2'h3;
    end else begin
      if (_T_3030) begin
        _T_3014 <= _T_3034;
      end
    end
    if (reset) begin
      _T_3107_0 <= 1'h0;
    end else begin
      if (_T_3003) begin
        _T_3107_0 <= _T_3046;
      end
    end
    if (reset) begin
      _T_3107_1 <= 1'h0;
    end else begin
      if (_T_3003) begin
        _T_3107_1 <= _T_3047;
      end
    end
    if (reset) begin
      _T_3180 <= 10'h0;
    end else begin
      if (_T_3183) begin
        _T_3180 <= _T_3285;
      end else begin
        _T_3180 <= _T_3289;
      end
    end
    if (reset) begin
      _T_3194 <= 3'h7;
    end else begin
      if (_T_3212) begin
        _T_3194 <= _T_3219;
      end
    end
    if (reset) begin
      _T_3312_0 <= 1'h0;
    end else begin
      if (_T_3182) begin
        _T_3312_0 <= _T_3233;
      end
    end
    if (reset) begin
      _T_3312_1 <= 1'h0;
    end else begin
      if (_T_3182) begin
        _T_3312_1 <= _T_3234;
      end
    end
    if (reset) begin
      _T_3312_2 <= 1'h0;
    end else begin
      if (_T_3182) begin
        _T_3312_2 <= _T_3235;
      end
    end
    if (reset) begin
      _T_3404 <= 10'h0;
    end else begin
      if (_T_3407) begin
        _T_3404 <= _T_3509;
      end else begin
        _T_3404 <= _T_3513;
      end
    end
    if (reset) begin
      _T_3418 <= 3'h7;
    end else begin
      if (_T_3436) begin
        _T_3418 <= _T_3443;
      end
    end
    if (reset) begin
      _T_3536_0 <= 1'h0;
    end else begin
      if (_T_3406) begin
        _T_3536_0 <= _T_3457;
      end
    end
    if (reset) begin
      _T_3536_1 <= 1'h0;
    end else begin
      if (_T_3406) begin
        _T_3536_1 <= _T_3458;
      end
    end
    if (reset) begin
      _T_3536_2 <= 1'h0;
    end else begin
      if (_T_3406) begin
        _T_3536_2 <= _T_3459;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2654) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2654) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2715) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2715) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2723) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2723) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2832) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2832) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2893) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2893) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2901) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2901) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3010) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3010) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3071) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3071) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3079) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3079) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3190) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3190) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3267) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3267) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3277) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3277) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3414) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3414) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3491) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3491) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3501) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3501) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [2:0] ram_param [0:0];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_35_data;
  wire  ram_param__T_35_addr;
  wire [2:0] ram_param__T_26_data;
  wire  ram_param__T_26_addr;
  wire  ram_param__T_26_mask;
  wire  ram_param__T_26_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_2;
  wire [2:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [2:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg [31:0] ram_address [0:0];
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_35_data;
  wire  ram_address__T_35_addr;
  wire [31:0] ram_address__T_26_data;
  wire  ram_address__T_26_addr;
  wire  ram_address__T_26_mask;
  wire  ram_address__T_26_en;
  reg [3:0] ram_mask [0:0];
  reg [31:0] _RAND_5;
  wire [3:0] ram_mask__T_35_data;
  wire  ram_mask__T_35_addr;
  wire [3:0] ram_mask__T_26_data;
  wire  ram_mask__T_26_addr;
  wire  ram_mask__T_26_mask;
  wire  ram_mask__T_26_en;
  reg [31:0] ram_data [0:0];
  reg [31:0] _RAND_6;
  wire [31:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [31:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  wire  _GEN_12;
  wire [2:0] _GEN_13;
  wire [2:0] _GEN_14;
  wire [2:0] _GEN_15;
  wire [4:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [3:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_11;
  assign io_deq_bits_opcode = _GEN_13;
  assign io_deq_bits_param = _GEN_14;
  assign io_deq_bits_size = _GEN_15;
  assign io_deq_bits_source = _GEN_16;
  assign io_deq_bits_address = _GEN_17;
  assign io_deq_bits_mask = _GEN_18;
  assign io_deq_bits_data = _GEN_19;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _GEN_21;
  assign ram_opcode__T_26_en = _GEN_21;
  assign ram_param__T_35_addr = 1'h0;
  assign ram_param__T_35_data = ram_param[ram_param__T_35_addr];
  assign ram_param__T_26_data = io_enq_bits_param;
  assign ram_param__T_26_addr = 1'h0;
  assign ram_param__T_26_mask = _GEN_21;
  assign ram_param__T_26_en = _GEN_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_21;
  assign ram_size__T_26_en = _GEN_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _GEN_21;
  assign ram_source__T_26_en = _GEN_21;
  assign ram_address__T_35_addr = 1'h0;
  assign ram_address__T_35_data = ram_address[ram_address__T_35_addr];
  assign ram_address__T_26_data = io_enq_bits_address;
  assign ram_address__T_26_addr = 1'h0;
  assign ram_address__T_26_mask = _GEN_21;
  assign ram_address__T_26_en = _GEN_21;
  assign ram_mask__T_35_addr = 1'h0;
  assign ram_mask__T_35_data = ram_mask[ram_mask__T_35_addr];
  assign ram_mask__T_26_data = io_enq_bits_mask;
  assign ram_mask__T_26_addr = 1'h0;
  assign ram_mask__T_26_mask = _GEN_21;
  assign ram_mask__T_26_en = _GEN_21;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _GEN_21;
  assign ram_data__T_26_en = _GEN_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_21 != _GEN_20;
  assign _GEN_10 = _T_29 ? _GEN_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_12 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_13 = _T_18 ? io_enq_bits_opcode : ram_opcode__T_35_data;
  assign _GEN_14 = _T_18 ? io_enq_bits_param : ram_param__T_35_data;
  assign _GEN_15 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_16 = _T_18 ? io_enq_bits_source : ram_source__T_35_data;
  assign _GEN_17 = _T_18 ? io_enq_bits_address : ram_address__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_mask : ram_mask__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_data : ram_data__T_35_data;
  assign _GEN_20 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_21 = _T_18 ? _GEN_12 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_param__T_26_en & ram_param__T_26_mask) begin
      ram_param[ram_param__T_26_addr] <= ram_param__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if(ram_address__T_26_en & ram_address__T_26_mask) begin
      ram_address[ram_address__T_26_addr] <= ram_address__T_26_data;
    end
    if(ram_mask__T_26_en & ram_mask__T_26_mask) begin
      ram_mask[ram_mask__T_26_addr] <= ram_mask__T_26_data;
    end
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input         io_enq_bits_sink,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output        io_deq_bits_sink,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [1:0] ram_param [0:0];
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_35_data;
  wire  ram_param__T_35_addr;
  wire [1:0] ram_param__T_26_data;
  wire  ram_param__T_26_addr;
  wire  ram_param__T_26_mask;
  wire  ram_param__T_26_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_2;
  wire [2:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [2:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  ram_sink [0:0];
  reg [31:0] _RAND_4;
  wire  ram_sink__T_35_data;
  wire  ram_sink__T_35_addr;
  wire  ram_sink__T_26_data;
  wire  ram_sink__T_26_addr;
  wire  ram_sink__T_26_mask;
  wire  ram_sink__T_26_en;
  reg [31:0] ram_data [0:0];
  reg [31:0] _RAND_5;
  wire [31:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [31:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg  ram_error [0:0];
  reg [31:0] _RAND_6;
  wire  ram_error__T_35_data;
  wire  ram_error__T_35_addr;
  wire  ram_error__T_26_data;
  wire  ram_error__T_26_addr;
  wire  ram_error__T_26_mask;
  wire  ram_error__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  wire  _GEN_12;
  wire [2:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [2:0] _GEN_15;
  wire [4:0] _GEN_16;
  wire  _GEN_17;
  wire [31:0] _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_11;
  assign io_deq_bits_opcode = _GEN_13;
  assign io_deq_bits_param = _GEN_14;
  assign io_deq_bits_size = _GEN_15;
  assign io_deq_bits_source = _GEN_16;
  assign io_deq_bits_sink = _GEN_17;
  assign io_deq_bits_data = _GEN_18;
  assign io_deq_bits_error = _GEN_19;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _GEN_21;
  assign ram_opcode__T_26_en = _GEN_21;
  assign ram_param__T_35_addr = 1'h0;
  assign ram_param__T_35_data = ram_param[ram_param__T_35_addr];
  assign ram_param__T_26_data = io_enq_bits_param;
  assign ram_param__T_26_addr = 1'h0;
  assign ram_param__T_26_mask = _GEN_21;
  assign ram_param__T_26_en = _GEN_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_21;
  assign ram_size__T_26_en = _GEN_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _GEN_21;
  assign ram_source__T_26_en = _GEN_21;
  assign ram_sink__T_35_addr = 1'h0;
  assign ram_sink__T_35_data = ram_sink[ram_sink__T_35_addr];
  assign ram_sink__T_26_data = io_enq_bits_sink;
  assign ram_sink__T_26_addr = 1'h0;
  assign ram_sink__T_26_mask = _GEN_21;
  assign ram_sink__T_26_en = _GEN_21;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _GEN_21;
  assign ram_data__T_26_en = _GEN_21;
  assign ram_error__T_35_addr = 1'h0;
  assign ram_error__T_35_data = ram_error[ram_error__T_35_addr];
  assign ram_error__T_26_data = io_enq_bits_error;
  assign ram_error__T_26_addr = 1'h0;
  assign ram_error__T_26_mask = _GEN_21;
  assign ram_error__T_26_en = _GEN_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_21 != _GEN_20;
  assign _GEN_10 = _T_29 ? _GEN_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_12 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_13 = _T_18 ? io_enq_bits_opcode : ram_opcode__T_35_data;
  assign _GEN_14 = _T_18 ? io_enq_bits_param : ram_param__T_35_data;
  assign _GEN_15 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_16 = _T_18 ? io_enq_bits_source : ram_source__T_35_data;
  assign _GEN_17 = _T_18 ? io_enq_bits_sink : ram_sink__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_data : ram_data__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_error : ram_error__T_35_data;
  assign _GEN_20 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_21 = _T_18 ? _GEN_12 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_error[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_param__T_26_en & ram_param__T_26_mask) begin
      ram_param[ram_param__T_26_addr] <= ram_param__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if(ram_sink__T_26_en & ram_sink__T_26_mask) begin
      ram_sink[ram_sink__T_26_addr] <= ram_sink__T_26_data;
    end
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if(ram_error__T_26_en & ram_error__T_26_mask) begin
      ram_error[ram_error__T_26_addr] <= ram_error__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [30:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [30:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_2;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg [30:0] ram_address [0:0];
  reg [31:0] _RAND_3;
  wire [30:0] ram_address__T_35_data;
  wire  ram_address__T_35_addr;
  wire [30:0] ram_address__T_26_data;
  wire  ram_address__T_26_addr;
  wire  ram_address__T_26_mask;
  wire  ram_address__T_26_en;
  reg [3:0] ram_mask [0:0];
  reg [31:0] _RAND_4;
  wire [3:0] ram_mask__T_35_data;
  wire  ram_mask__T_35_addr;
  wire [3:0] ram_mask__T_26_data;
  wire  ram_mask__T_26_addr;
  wire  ram_mask__T_26_mask;
  wire  ram_mask__T_26_en;
  reg [31:0] ram_data [0:0];
  reg [31:0] _RAND_5;
  wire [31:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [31:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_6;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  wire  _GEN_12;
  wire [2:0] _GEN_13;
  wire [3:0] _GEN_15;
  wire [4:0] _GEN_16;
  wire [30:0] _GEN_17;
  wire [3:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_11;
  assign io_deq_bits_opcode = _GEN_13;
  assign io_deq_bits_size = _GEN_15;
  assign io_deq_bits_source = _GEN_16;
  assign io_deq_bits_address = _GEN_17;
  assign io_deq_bits_mask = _GEN_18;
  assign io_deq_bits_data = _GEN_19;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _GEN_21;
  assign ram_opcode__T_26_en = _GEN_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_21;
  assign ram_size__T_26_en = _GEN_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _GEN_21;
  assign ram_source__T_26_en = _GEN_21;
  assign ram_address__T_35_addr = 1'h0;
  assign ram_address__T_35_data = ram_address[ram_address__T_35_addr];
  assign ram_address__T_26_data = io_enq_bits_address;
  assign ram_address__T_26_addr = 1'h0;
  assign ram_address__T_26_mask = _GEN_21;
  assign ram_address__T_26_en = _GEN_21;
  assign ram_mask__T_35_addr = 1'h0;
  assign ram_mask__T_35_data = ram_mask[ram_mask__T_35_addr];
  assign ram_mask__T_26_data = io_enq_bits_mask;
  assign ram_mask__T_26_addr = 1'h0;
  assign ram_mask__T_26_mask = _GEN_21;
  assign ram_mask__T_26_en = _GEN_21;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _GEN_21;
  assign ram_data__T_26_en = _GEN_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_21 != _GEN_20;
  assign _GEN_10 = _T_29 ? _GEN_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_12 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_13 = _T_18 ? io_enq_bits_opcode : ram_opcode__T_35_data;
  assign _GEN_15 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_16 = _T_18 ? io_enq_bits_source : ram_source__T_35_data;
  assign _GEN_17 = _T_18 ? io_enq_bits_address : ram_address__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_mask : ram_mask__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_data : ram_data__T_35_data;
  assign _GEN_20 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_21 = _T_18 ? _GEN_12 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_address[initvar] = _RAND_3[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask[initvar] = _RAND_4[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  maybe_full = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if(ram_address__T_26_en & ram_address__T_26_mask) begin
      ram_address[ram_address__T_26_addr] <= ram_address__T_26_data;
    end
    if(ram_mask__T_26_en & ram_mask__T_26_mask) begin
      ram_mask[ram_mask__T_26_addr] <= ram_mask__T_26_data;
    end
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input         io_enq_bits_sink,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output        io_deq_bits_sink,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [1:0] ram_param [0:0];
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_35_data;
  wire  ram_param__T_35_addr;
  wire [1:0] ram_param__T_26_data;
  wire  ram_param__T_26_addr;
  wire  ram_param__T_26_mask;
  wire  ram_param__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  ram_sink [0:0];
  reg [31:0] _RAND_4;
  wire  ram_sink__T_35_data;
  wire  ram_sink__T_35_addr;
  wire  ram_sink__T_26_data;
  wire  ram_sink__T_26_addr;
  wire  ram_sink__T_26_mask;
  wire  ram_sink__T_26_en;
  reg [31:0] ram_data [0:0];
  reg [31:0] _RAND_5;
  wire [31:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [31:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg  ram_error [0:0];
  reg [31:0] _RAND_6;
  wire  ram_error__T_35_data;
  wire  ram_error__T_35_addr;
  wire  ram_error__T_26_data;
  wire  ram_error__T_26_addr;
  wire  ram_error__T_26_mask;
  wire  ram_error__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  wire  _GEN_12;
  wire [2:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [3:0] _GEN_15;
  wire [4:0] _GEN_16;
  wire  _GEN_17;
  wire [31:0] _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_11;
  assign io_deq_bits_opcode = _GEN_13;
  assign io_deq_bits_param = _GEN_14;
  assign io_deq_bits_size = _GEN_15;
  assign io_deq_bits_source = _GEN_16;
  assign io_deq_bits_sink = _GEN_17;
  assign io_deq_bits_data = _GEN_18;
  assign io_deq_bits_error = _GEN_19;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _GEN_21;
  assign ram_opcode__T_26_en = _GEN_21;
  assign ram_param__T_35_addr = 1'h0;
  assign ram_param__T_35_data = ram_param[ram_param__T_35_addr];
  assign ram_param__T_26_data = io_enq_bits_param;
  assign ram_param__T_26_addr = 1'h0;
  assign ram_param__T_26_mask = _GEN_21;
  assign ram_param__T_26_en = _GEN_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_21;
  assign ram_size__T_26_en = _GEN_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _GEN_21;
  assign ram_source__T_26_en = _GEN_21;
  assign ram_sink__T_35_addr = 1'h0;
  assign ram_sink__T_35_data = ram_sink[ram_sink__T_35_addr];
  assign ram_sink__T_26_data = io_enq_bits_sink;
  assign ram_sink__T_26_addr = 1'h0;
  assign ram_sink__T_26_mask = _GEN_21;
  assign ram_sink__T_26_en = _GEN_21;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _GEN_21;
  assign ram_data__T_26_en = _GEN_21;
  assign ram_error__T_35_addr = 1'h0;
  assign ram_error__T_35_data = ram_error[ram_error__T_35_addr];
  assign ram_error__T_26_data = io_enq_bits_error;
  assign ram_error__T_26_addr = 1'h0;
  assign ram_error__T_26_mask = _GEN_21;
  assign ram_error__T_26_en = _GEN_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_21 != _GEN_20;
  assign _GEN_10 = _T_29 ? _GEN_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_12 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_13 = _T_18 ? io_enq_bits_opcode : ram_opcode__T_35_data;
  assign _GEN_14 = _T_18 ? io_enq_bits_param : ram_param__T_35_data;
  assign _GEN_15 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_16 = _T_18 ? io_enq_bits_source : ram_source__T_35_data;
  assign _GEN_17 = _T_18 ? io_enq_bits_sink : ram_sink__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_data : ram_data__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_error : ram_error__T_35_data;
  assign _GEN_20 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_21 = _T_18 ? _GEN_12 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_error[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_param__T_26_en & ram_param__T_26_mask) begin
      ram_param[ram_param__T_26_addr] <= ram_param__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if(ram_sink__T_26_en & ram_sink__T_26_mask) begin
      ram_sink[ram_sink__T_26_addr] <= ram_sink__T_26_data;
    end
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if(ram_error__T_26_en & ram_error__T_26_mask) begin
      ram_error[ram_error__T_26_addr] <= ram_error__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_4(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [3:0] io_enq_bits_size,
  input  [4:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_2;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  wire  _GEN_12;
  wire [2:0] _GEN_13;
  wire [3:0] _GEN_15;
  wire [4:0] _GEN_16;
  wire  _GEN_20;
  wire  _GEN_21;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_11;
  assign io_deq_bits_opcode = _GEN_13;
  assign io_deq_bits_size = _GEN_15;
  assign io_deq_bits_source = _GEN_16;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _GEN_21;
  assign ram_opcode__T_26_en = _GEN_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_21;
  assign ram_size__T_26_en = _GEN_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _GEN_21;
  assign ram_source__T_26_en = _GEN_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_21 != _GEN_20;
  assign _GEN_10 = _T_29 ? _GEN_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_12 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_13 = _T_18 ? io_enq_bits_opcode : ram_opcode__T_35_data;
  assign _GEN_15 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_16 = _T_18 ? io_enq_bits_source : ram_source__T_35_data;
  assign _GEN_20 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_21 = _T_18 ? _GEN_12 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module TLBuffer_1(
  input         clock,
  input         reset,
  output        io_in_2_a_ready,
  input         io_in_2_a_valid,
  input  [2:0]  io_in_2_a_bits_opcode,
  input  [3:0]  io_in_2_a_bits_size,
  input  [4:0]  io_in_2_a_bits_source,
  input         io_in_2_d_ready,
  output        io_in_2_d_valid,
  output [2:0]  io_in_2_d_bits_opcode,
  output [1:0]  io_in_2_d_bits_param,
  output [3:0]  io_in_2_d_bits_size,
  output [4:0]  io_in_2_d_bits_source,
  output        io_in_2_d_bits_sink,
  output [31:0] io_in_2_d_bits_data,
  output        io_in_2_d_bits_error,
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [3:0]  io_in_1_a_bits_size,
  input  [4:0]  io_in_1_a_bits_source,
  input  [30:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [1:0]  io_in_1_d_bits_param,
  output [3:0]  io_in_1_d_bits_size,
  output [4:0]  io_in_1_d_bits_source,
  output        io_in_1_d_bits_sink,
  output [31:0] io_in_1_d_bits_data,
  output        io_in_1_d_bits_error,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_2_a_ready,
  output        io_out_2_a_valid,
  output [2:0]  io_out_2_a_bits_opcode,
  output [3:0]  io_out_2_a_bits_size,
  output [4:0]  io_out_2_a_bits_source,
  output        io_out_2_d_ready,
  input         io_out_2_d_valid,
  input  [2:0]  io_out_2_d_bits_opcode,
  input  [1:0]  io_out_2_d_bits_param,
  input  [3:0]  io_out_2_d_bits_size,
  input  [4:0]  io_out_2_d_bits_source,
  input         io_out_2_d_bits_sink,
  input  [31:0] io_out_2_d_bits_data,
  input         io_out_2_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [3:0]  io_out_1_a_bits_size,
  output [4:0]  io_out_1_a_bits_source,
  output [30:0] io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [3:0]  io_out_1_d_bits_size,
  input  [4:0]  io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [31:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [2:0] Queue_io_enq_bits_param;
  wire [2:0] Queue_io_enq_bits_size;
  wire [4:0] Queue_io_enq_bits_source;
  wire [31:0] Queue_io_enq_bits_address;
  wire [3:0] Queue_io_enq_bits_mask;
  wire [31:0] Queue_io_enq_bits_data;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [2:0] Queue_io_deq_bits_param;
  wire [2:0] Queue_io_deq_bits_size;
  wire [4:0] Queue_io_deq_bits_source;
  wire [31:0] Queue_io_deq_bits_address;
  wire [3:0] Queue_io_deq_bits_mask;
  wire [31:0] Queue_io_deq_bits_data;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [1:0] Queue_1_io_enq_bits_param;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [4:0] Queue_1_io_enq_bits_source;
  wire  Queue_1_io_enq_bits_sink;
  wire [31:0] Queue_1_io_enq_bits_data;
  wire  Queue_1_io_enq_bits_error;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [1:0] Queue_1_io_deq_bits_param;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [4:0] Queue_1_io_deq_bits_source;
  wire  Queue_1_io_deq_bits_sink;
  wire [31:0] Queue_1_io_deq_bits_data;
  wire  Queue_1_io_deq_bits_error;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [2:0] Queue_2_io_enq_bits_opcode;
  wire [3:0] Queue_2_io_enq_bits_size;
  wire [4:0] Queue_2_io_enq_bits_source;
  wire [30:0] Queue_2_io_enq_bits_address;
  wire [3:0] Queue_2_io_enq_bits_mask;
  wire [31:0] Queue_2_io_enq_bits_data;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [2:0] Queue_2_io_deq_bits_opcode;
  wire [3:0] Queue_2_io_deq_bits_size;
  wire [4:0] Queue_2_io_deq_bits_source;
  wire [30:0] Queue_2_io_deq_bits_address;
  wire [3:0] Queue_2_io_deq_bits_mask;
  wire [31:0] Queue_2_io_deq_bits_data;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [2:0] Queue_3_io_enq_bits_opcode;
  wire [1:0] Queue_3_io_enq_bits_param;
  wire [3:0] Queue_3_io_enq_bits_size;
  wire [4:0] Queue_3_io_enq_bits_source;
  wire  Queue_3_io_enq_bits_sink;
  wire [31:0] Queue_3_io_enq_bits_data;
  wire  Queue_3_io_enq_bits_error;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [2:0] Queue_3_io_deq_bits_opcode;
  wire [1:0] Queue_3_io_deq_bits_param;
  wire [3:0] Queue_3_io_deq_bits_size;
  wire [4:0] Queue_3_io_deq_bits_source;
  wire  Queue_3_io_deq_bits_sink;
  wire [31:0] Queue_3_io_deq_bits_data;
  wire  Queue_3_io_deq_bits_error;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [2:0] Queue_4_io_enq_bits_opcode;
  wire [3:0] Queue_4_io_enq_bits_size;
  wire [4:0] Queue_4_io_enq_bits_source;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [2:0] Queue_4_io_deq_bits_opcode;
  wire [3:0] Queue_4_io_deq_bits_size;
  wire [4:0] Queue_4_io_deq_bits_source;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire [2:0] Queue_5_io_enq_bits_opcode;
  wire [1:0] Queue_5_io_enq_bits_param;
  wire [3:0] Queue_5_io_enq_bits_size;
  wire [4:0] Queue_5_io_enq_bits_source;
  wire  Queue_5_io_enq_bits_sink;
  wire [31:0] Queue_5_io_enq_bits_data;
  wire  Queue_5_io_enq_bits_error;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire [2:0] Queue_5_io_deq_bits_opcode;
  wire [1:0] Queue_5_io_deq_bits_param;
  wire [3:0] Queue_5_io_deq_bits_size;
  wire [4:0] Queue_5_io_deq_bits_source;
  wire  Queue_5_io_deq_bits_sink;
  wire [31:0] Queue_5_io_deq_bits_data;
  wire  Queue_5_io_deq_bits_error;
  Queue Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_1 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_error(Queue_1_io_enq_bits_error),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_error(Queue_1_io_deq_bits_error)
  );
  Queue_2 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_opcode(Queue_2_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_2_io_enq_bits_size),
    .io_enq_bits_source(Queue_2_io_enq_bits_source),
    .io_enq_bits_address(Queue_2_io_enq_bits_address),
    .io_enq_bits_mask(Queue_2_io_enq_bits_mask),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_opcode(Queue_2_io_deq_bits_opcode),
    .io_deq_bits_size(Queue_2_io_deq_bits_size),
    .io_deq_bits_source(Queue_2_io_deq_bits_source),
    .io_deq_bits_address(Queue_2_io_deq_bits_address),
    .io_deq_bits_mask(Queue_2_io_deq_bits_mask),
    .io_deq_bits_data(Queue_2_io_deq_bits_data)
  );
  Queue_3 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_opcode(Queue_3_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_3_io_enq_bits_param),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_source(Queue_3_io_enq_bits_source),
    .io_enq_bits_sink(Queue_3_io_enq_bits_sink),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_enq_bits_error(Queue_3_io_enq_bits_error),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_opcode(Queue_3_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_3_io_deq_bits_param),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_source(Queue_3_io_deq_bits_source),
    .io_deq_bits_sink(Queue_3_io_deq_bits_sink),
    .io_deq_bits_data(Queue_3_io_deq_bits_data),
    .io_deq_bits_error(Queue_3_io_deq_bits_error)
  );
  Queue_4 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_opcode(Queue_4_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_4_io_enq_bits_size),
    .io_enq_bits_source(Queue_4_io_enq_bits_source),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_opcode(Queue_4_io_deq_bits_opcode),
    .io_deq_bits_size(Queue_4_io_deq_bits_size),
    .io_deq_bits_source(Queue_4_io_deq_bits_source)
  );
  Queue_3 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits_opcode(Queue_5_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_5_io_enq_bits_param),
    .io_enq_bits_size(Queue_5_io_enq_bits_size),
    .io_enq_bits_source(Queue_5_io_enq_bits_source),
    .io_enq_bits_sink(Queue_5_io_enq_bits_sink),
    .io_enq_bits_data(Queue_5_io_enq_bits_data),
    .io_enq_bits_error(Queue_5_io_enq_bits_error),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits_opcode(Queue_5_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_5_io_deq_bits_param),
    .io_deq_bits_size(Queue_5_io_deq_bits_size),
    .io_deq_bits_source(Queue_5_io_deq_bits_source),
    .io_deq_bits_sink(Queue_5_io_deq_bits_sink),
    .io_deq_bits_data(Queue_5_io_deq_bits_data),
    .io_deq_bits_error(Queue_5_io_deq_bits_error)
  );
  assign io_in_2_a_ready = Queue_4_io_enq_ready;
  assign io_in_2_d_valid = Queue_5_io_deq_valid;
  assign io_in_2_d_bits_opcode = Queue_5_io_deq_bits_opcode;
  assign io_in_2_d_bits_param = Queue_5_io_deq_bits_param;
  assign io_in_2_d_bits_size = Queue_5_io_deq_bits_size;
  assign io_in_2_d_bits_source = Queue_5_io_deq_bits_source;
  assign io_in_2_d_bits_sink = Queue_5_io_deq_bits_sink;
  assign io_in_2_d_bits_data = Queue_5_io_deq_bits_data;
  assign io_in_2_d_bits_error = Queue_5_io_deq_bits_error;
  assign io_in_1_a_ready = Queue_2_io_enq_ready;
  assign io_in_1_d_valid = Queue_3_io_deq_valid;
  assign io_in_1_d_bits_opcode = Queue_3_io_deq_bits_opcode;
  assign io_in_1_d_bits_param = Queue_3_io_deq_bits_param;
  assign io_in_1_d_bits_size = Queue_3_io_deq_bits_size;
  assign io_in_1_d_bits_source = Queue_3_io_deq_bits_source;
  assign io_in_1_d_bits_sink = Queue_3_io_deq_bits_sink;
  assign io_in_1_d_bits_data = Queue_3_io_deq_bits_data;
  assign io_in_1_d_bits_error = Queue_3_io_deq_bits_error;
  assign io_in_0_a_ready = Queue_io_enq_ready;
  assign io_in_0_d_valid = Queue_1_io_deq_valid;
  assign io_in_0_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign io_in_0_d_bits_param = Queue_1_io_deq_bits_param;
  assign io_in_0_d_bits_size = Queue_1_io_deq_bits_size;
  assign io_in_0_d_bits_source = Queue_1_io_deq_bits_source;
  assign io_in_0_d_bits_sink = Queue_1_io_deq_bits_sink;
  assign io_in_0_d_bits_data = Queue_1_io_deq_bits_data;
  assign io_in_0_d_bits_error = Queue_1_io_deq_bits_error;
  assign io_out_2_a_valid = Queue_4_io_deq_valid;
  assign io_out_2_a_bits_opcode = Queue_4_io_deq_bits_opcode;
  assign io_out_2_a_bits_size = Queue_4_io_deq_bits_size;
  assign io_out_2_a_bits_source = Queue_4_io_deq_bits_source;
  assign io_out_2_d_ready = Queue_5_io_enq_ready;
  assign io_out_1_a_valid = Queue_2_io_deq_valid;
  assign io_out_1_a_bits_opcode = Queue_2_io_deq_bits_opcode;
  assign io_out_1_a_bits_size = Queue_2_io_deq_bits_size;
  assign io_out_1_a_bits_source = Queue_2_io_deq_bits_source;
  assign io_out_1_a_bits_address = Queue_2_io_deq_bits_address;
  assign io_out_1_a_bits_mask = Queue_2_io_deq_bits_mask;
  assign io_out_1_a_bits_data = Queue_2_io_deq_bits_data;
  assign io_out_1_d_ready = Queue_3_io_enq_ready;
  assign io_out_0_a_valid = Queue_io_deq_valid;
  assign io_out_0_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign io_out_0_a_bits_param = Queue_io_deq_bits_param;
  assign io_out_0_a_bits_size = Queue_io_deq_bits_size;
  assign io_out_0_a_bits_source = Queue_io_deq_bits_source;
  assign io_out_0_a_bits_address = Queue_io_deq_bits_address;
  assign io_out_0_a_bits_mask = Queue_io_deq_bits_mask;
  assign io_out_0_a_bits_data = Queue_io_deq_bits_data;
  assign io_out_0_d_ready = Queue_1_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_a_valid;
  assign Queue_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Queue_io_enq_bits_param = io_in_0_a_bits_param;
  assign Queue_io_enq_bits_size = io_in_0_a_bits_size;
  assign Queue_io_enq_bits_source = io_in_0_a_bits_source;
  assign Queue_io_enq_bits_address = io_in_0_a_bits_address;
  assign Queue_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Queue_io_enq_bits_data = io_in_0_a_bits_data;
  assign Queue_io_deq_ready = io_out_0_a_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_out_0_d_valid;
  assign Queue_1_io_enq_bits_opcode = io_out_0_d_bits_opcode;
  assign Queue_1_io_enq_bits_param = io_out_0_d_bits_param;
  assign Queue_1_io_enq_bits_size = io_out_0_d_bits_size;
  assign Queue_1_io_enq_bits_source = io_out_0_d_bits_source;
  assign Queue_1_io_enq_bits_sink = io_out_0_d_bits_sink;
  assign Queue_1_io_enq_bits_data = io_out_0_d_bits_data;
  assign Queue_1_io_enq_bits_error = io_out_0_d_bits_error;
  assign Queue_1_io_deq_ready = io_in_0_d_ready;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = io_in_1_a_valid;
  assign Queue_2_io_enq_bits_opcode = io_in_1_a_bits_opcode;
  assign Queue_2_io_enq_bits_size = io_in_1_a_bits_size;
  assign Queue_2_io_enq_bits_source = io_in_1_a_bits_source;
  assign Queue_2_io_enq_bits_address = io_in_1_a_bits_address;
  assign Queue_2_io_enq_bits_mask = io_in_1_a_bits_mask;
  assign Queue_2_io_enq_bits_data = io_in_1_a_bits_data;
  assign Queue_2_io_deq_ready = io_out_1_a_ready;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = io_out_1_d_valid;
  assign Queue_3_io_enq_bits_opcode = io_out_1_d_bits_opcode;
  assign Queue_3_io_enq_bits_param = io_out_1_d_bits_param;
  assign Queue_3_io_enq_bits_size = io_out_1_d_bits_size;
  assign Queue_3_io_enq_bits_source = io_out_1_d_bits_source;
  assign Queue_3_io_enq_bits_sink = io_out_1_d_bits_sink;
  assign Queue_3_io_enq_bits_data = io_out_1_d_bits_data;
  assign Queue_3_io_enq_bits_error = io_out_1_d_bits_error;
  assign Queue_3_io_deq_ready = io_in_1_d_ready;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = io_in_2_a_valid;
  assign Queue_4_io_enq_bits_opcode = io_in_2_a_bits_opcode;
  assign Queue_4_io_enq_bits_size = io_in_2_a_bits_size;
  assign Queue_4_io_enq_bits_source = io_in_2_a_bits_source;
  assign Queue_4_io_deq_ready = io_out_2_a_ready;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_5_io_enq_valid = io_out_2_d_valid;
  assign Queue_5_io_enq_bits_opcode = io_out_2_d_bits_opcode;
  assign Queue_5_io_enq_bits_param = io_out_2_d_bits_param;
  assign Queue_5_io_enq_bits_size = io_out_2_d_bits_size;
  assign Queue_5_io_enq_bits_source = io_out_2_d_bits_source;
  assign Queue_5_io_enq_bits_sink = io_out_2_d_bits_sink;
  assign Queue_5_io_enq_bits_data = io_out_2_d_bits_data;
  assign Queue_5_io_enq_bits_error = io_out_2_d_bits_error;
  assign Queue_5_io_deq_ready = io_in_2_d_ready;
endmodule
module Repeater(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input         io_enq_bits_sink,
  input  [63:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output        io_deq_bits_sink,
  output [63:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [1:0] saved_param;
  reg [31:0] _RAND_2;
  reg [3:0] saved_size;
  reg [31:0] _RAND_3;
  reg [4:0] saved_source;
  reg [31:0] _RAND_4;
  reg  saved_sink;
  reg [31:0] _RAND_5;
  reg [63:0] saved_data;
  reg [63:0] _RAND_6;
  reg  saved_error;
  reg [31:0] _RAND_7;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [1:0] _T_20_param;
  wire [3:0] _T_20_size;
  wire [4:0] _T_20_source;
  wire  _T_20_sink;
  wire [63:0] _T_20_data;
  wire  _T_20_error;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [1:0] _GEN_2;
  wire [3:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire  _GEN_5;
  wire [63:0] _GEN_6;
  wire  _GEN_7;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_param = _T_20_param;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_sink = _T_20_sink;
  assign io_deq_bits_data = _T_20_data;
  assign io_deq_bits_error = _T_20_error;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_param = full ? saved_param : io_enq_bits_param;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_sink = full ? saved_sink : io_enq_bits_sink;
  assign _T_20_data = full ? saved_data : io_enq_bits_data;
  assign _T_20_error = full ? saved_error : io_enq_bits_error;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_2 = _T_22 ? io_enq_bits_param : saved_param;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_sink : saved_sink;
  assign _GEN_6 = _T_22 ? io_enq_bits_data : saved_data;
  assign _GEN_7 = _T_22 ? io_enq_bits_error : saved_error;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_param = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_size = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_source = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_sink = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{$random}};
  saved_data = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  saved_error = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_sink <= io_enq_bits_sink;
    end
    if (_T_22) begin
      saved_data <= io_enq_bits_data;
    end
    if (_T_22) begin
      saved_error <= io_enq_bits_error;
    end
  end
endmodule
module TLWidthWidget(
  input         clock,
  input         reset,
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [3:0]  io_in_1_a_bits_size,
  input  [4:0]  io_in_1_a_bits_source,
  input  [30:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [1:0]  io_in_1_d_bits_param,
  output [3:0]  io_in_1_d_bits_size,
  output [4:0]  io_in_1_d_bits_source,
  output        io_in_1_d_bits_sink,
  output [31:0] io_in_1_d_bits_data,
  output        io_in_1_d_bits_error,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [3:0]  io_out_1_a_bits_size,
  output [4:0]  io_out_1_a_bits_source,
  output [30:0] io_out_1_a_bits_address,
  output [7:0]  io_out_1_a_bits_mask,
  output [63:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [3:0]  io_out_1_d_bits_size,
  input  [4:0]  io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [63:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  _T_183;
  wire  _T_185;
  wire [17:0] _T_188;
  wire [2:0] _T_189;
  wire [2:0] _T_190;
  wire  _T_191;
  reg  _T_194;
  reg [31:0] _RAND_0;
  wire  _T_197;
  wire  _T_199;
  wire  _T_200;
  wire  _T_203;
  wire  _T_207;
  wire  _T_215;
  wire [1:0] _T_217;
  wire  _T_218;
  wire  _GEN_3;
  wire  _GEN_4;
  wire  _T_221;
  wire  _T_222;
  wire  _T_223;
  reg [31:0] _T_226_0;
  reg [31:0] _RAND_1;
  wire [31:0] _T_230;
  wire  _T_235;
  wire [31:0] _GEN_5;
  wire [63:0] _T_236;
  wire [1:0] _T_237;
  wire [3:0] _T_239;
  wire [2:0] _T_240;
  wire [2:0] _T_242;
  wire  _T_244;
  wire  _T_246;
  wire  _T_247;
  wire  _T_249;
  wire  _T_251;
  wire  _T_252;
  wire  _T_254;
  wire  _T_255;
  wire  _T_256;
  wire  _T_257;
  wire  _T_259;
  wire  _T_260;
  wire  _T_261;
  wire  _T_262;
  wire  _T_263;
  wire  _T_264;
  wire  _T_265;
  wire  _T_266;
  wire  _T_267;
  wire  _T_268;
  wire  _T_269;
  wire  _T_270;
  wire  _T_271;
  wire  _T_272;
  wire  _T_273;
  wire  _T_275;
  wire  _T_276;
  wire  _T_277;
  wire  _T_278;
  wire  _T_279;
  wire  _T_280;
  wire  _T_281;
  wire  _T_282;
  wire  _T_283;
  wire  _T_284;
  wire  _T_285;
  wire  _T_286;
  wire  _T_287;
  wire  _T_288;
  wire  _T_289;
  wire  _T_290;
  wire  _T_291;
  wire  _T_292;
  wire  _T_293;
  wire  _T_294;
  wire  _T_295;
  wire  _T_296;
  wire  _T_297;
  wire  _T_298;
  wire  _T_299;
  wire [1:0] _T_300;
  wire [1:0] _T_301;
  wire [3:0] _T_302;
  wire [1:0] _T_303;
  wire [1:0] _T_304;
  wire [3:0] _T_305;
  wire [7:0] _T_306;
  reg [3:0] _T_309_0;
  reg [31:0] _RAND_2;
  wire [3:0] _T_313;
  wire [3:0] _GEN_6;
  wire [7:0] _T_319;
  wire [7:0] _T_322;
  wire [7:0] _T_323;
  wire  Repeater_clock;
  wire  Repeater_reset;
  wire  Repeater_io_repeat;
  wire  Repeater_io_enq_ready;
  wire  Repeater_io_enq_valid;
  wire [2:0] Repeater_io_enq_bits_opcode;
  wire [1:0] Repeater_io_enq_bits_param;
  wire [3:0] Repeater_io_enq_bits_size;
  wire [4:0] Repeater_io_enq_bits_source;
  wire  Repeater_io_enq_bits_sink;
  wire [63:0] Repeater_io_enq_bits_data;
  wire  Repeater_io_enq_bits_error;
  wire  Repeater_io_deq_ready;
  wire  Repeater_io_deq_valid;
  wire [2:0] Repeater_io_deq_bits_opcode;
  wire [1:0] Repeater_io_deq_bits_param;
  wire [3:0] Repeater_io_deq_bits_size;
  wire [4:0] Repeater_io_deq_bits_source;
  wire  Repeater_io_deq_bits_sink;
  wire [63:0] Repeater_io_deq_bits_data;
  wire  Repeater_io_deq_bits_error;
  wire  _T_326_valid;
  wire [2:0] _T_326_bits_opcode;
  wire [1:0] _T_326_bits_param;
  wire [3:0] _T_326_bits_size;
  wire [4:0] _T_326_bits_source;
  wire  _T_326_bits_sink;
  wire  _T_326_bits_error;
  wire [31:0] _T_330;
  wire [31:0] _T_331;
  wire [63:0] _T_332;
  wire  _T_333;
  wire [17:0] _T_336;
  wire [2:0] _T_337;
  wire [2:0] _T_338;
  wire  _T_339;
  reg  _T_342;
  reg [31:0] _RAND_3;
  wire  _T_344;
  wire  _T_345;
  wire  _T_347;
  wire  _T_348;
  wire  _T_349;
  wire [1:0] _T_351;
  wire  _T_352;
  wire  _GEN_7;
  wire  _GEN_8;
  reg  _T_357_0;
  reg [31:0] _RAND_4;
  reg  _T_357_1;
  reg [31:0] _RAND_5;
  reg  _T_357_2;
  reg [31:0] _RAND_6;
  reg  _T_357_3;
  reg [31:0] _RAND_7;
  reg  _T_357_4;
  reg [31:0] _RAND_8;
  reg  _T_357_5;
  reg [31:0] _RAND_9;
  reg  _T_357_6;
  reg [31:0] _RAND_10;
  reg  _T_357_7;
  reg [31:0] _RAND_11;
  reg  _T_357_8;
  reg [31:0] _RAND_12;
  reg  _T_357_9;
  reg [31:0] _RAND_13;
  reg  _T_357_10;
  reg [31:0] _RAND_14;
  reg  _T_357_11;
  reg [31:0] _RAND_15;
  reg  _T_357_12;
  reg [31:0] _RAND_16;
  reg  _T_357_13;
  reg [31:0] _RAND_17;
  reg  _T_357_14;
  reg [31:0] _RAND_18;
  reg  _T_357_15;
  reg [31:0] _RAND_19;
  reg  _T_357_16;
  reg [31:0] _RAND_20;
  reg  _T_357_17;
  reg [31:0] _RAND_21;
  wire  _T_378;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  reg  _T_389;
  reg [31:0] _RAND_22;
  wire  _GEN_62;
  wire  _T_391;
  wire  _T_392;
  wire  _T_393;
  wire [31:0] _T_394;
  wire [31:0] _T_395;
  wire [31:0] _GEN_63;
  wire  _T_405;
  Repeater Repeater (
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_io_enq_bits_param),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_sink(Repeater_io_enq_bits_sink),
    .io_enq_bits_data(Repeater_io_enq_bits_data),
    .io_enq_bits_error(Repeater_io_enq_bits_error),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_io_deq_bits_param),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_sink(Repeater_io_deq_bits_sink),
    .io_deq_bits_data(Repeater_io_deq_bits_data),
    .io_deq_bits_error(Repeater_io_deq_bits_error)
  );
  assign io_in_1_a_ready = _T_222;
  assign io_in_1_d_valid = _T_326_valid;
  assign io_in_1_d_bits_opcode = _T_326_bits_opcode;
  assign io_in_1_d_bits_param = _T_326_bits_param;
  assign io_in_1_d_bits_size = _T_326_bits_size;
  assign io_in_1_d_bits_source = _T_326_bits_source;
  assign io_in_1_d_bits_sink = _T_326_bits_sink;
  assign io_in_1_d_bits_data = _GEN_63;
  assign io_in_1_d_bits_error = _T_326_bits_error;
  assign io_in_0_a_ready = io_out_0_a_ready;
  assign io_in_0_d_valid = io_out_0_d_valid;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_param = io_out_0_d_bits_param;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_in_0_d_bits_sink = io_out_0_d_bits_sink;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_d_bits_error = io_out_0_d_bits_error;
  assign io_out_1_a_valid = _T_223;
  assign io_out_1_a_bits_opcode = io_in_1_a_bits_opcode;
  assign io_out_1_a_bits_size = io_in_1_a_bits_size;
  assign io_out_1_a_bits_source = io_in_1_a_bits_source;
  assign io_out_1_a_bits_address = io_in_1_a_bits_address;
  assign io_out_1_a_bits_mask = _T_323;
  assign io_out_1_a_bits_data = _T_236;
  assign io_out_1_d_ready = Repeater_io_enq_ready;
  assign io_out_0_a_valid = io_in_0_a_valid;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_param = io_in_0_a_bits_param;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address;
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = io_in_0_d_ready;
  assign _T_183 = io_in_1_a_bits_opcode[2];
  assign _T_185 = _T_183 == 1'h0;
  assign _T_188 = 18'h7 << io_in_1_a_bits_size;
  assign _T_189 = _T_188[2:0];
  assign _T_190 = ~ _T_189;
  assign _T_191 = _T_190[2:2];
  assign _T_197 = _T_194 == _T_191;
  assign _T_199 = _T_185 == 1'h0;
  assign _T_200 = _T_197 | _T_199;
  assign _T_203 = _T_194 & _T_191;
  assign _T_207 = _T_203 == 1'h0;
  assign _T_215 = io_in_1_a_ready & io_in_1_a_valid;
  assign _T_217 = _T_194 + 1'h1;
  assign _T_218 = _T_217[0:0];
  assign _GEN_3 = _T_200 ? 1'h0 : _T_218;
  assign _GEN_4 = _T_215 ? _GEN_3 : _T_194;
  assign _T_221 = _T_200 == 1'h0;
  assign _T_222 = io_out_1_a_ready | _T_221;
  assign _T_223 = io_in_1_a_valid & _T_200;
  assign _T_230 = _T_207 ? io_in_1_a_bits_data : _T_226_0;
  assign _T_235 = _T_215 & _T_221;
  assign _GEN_5 = _T_235 ? _T_230 : _T_226_0;
  assign _T_236 = {io_in_1_a_bits_data,_T_230};
  assign _T_237 = io_out_1_a_bits_size[1:0];
  assign _T_239 = 4'h1 << _T_237;
  assign _T_240 = _T_239[2:0];
  assign _T_242 = _T_240 | 3'h1;
  assign _T_244 = io_out_1_a_bits_size >= 4'h3;
  assign _T_246 = _T_242[2];
  assign _T_247 = io_out_1_a_bits_address[2];
  assign _T_249 = _T_247 == 1'h0;
  assign _T_251 = _T_246 & _T_249;
  assign _T_252 = _T_244 | _T_251;
  assign _T_254 = _T_246 & _T_247;
  assign _T_255 = _T_244 | _T_254;
  assign _T_256 = _T_242[1];
  assign _T_257 = io_out_1_a_bits_address[1];
  assign _T_259 = _T_257 == 1'h0;
  assign _T_260 = _T_249 & _T_259;
  assign _T_261 = _T_256 & _T_260;
  assign _T_262 = _T_252 | _T_261;
  assign _T_263 = _T_249 & _T_257;
  assign _T_264 = _T_256 & _T_263;
  assign _T_265 = _T_252 | _T_264;
  assign _T_266 = _T_247 & _T_259;
  assign _T_267 = _T_256 & _T_266;
  assign _T_268 = _T_255 | _T_267;
  assign _T_269 = _T_247 & _T_257;
  assign _T_270 = _T_256 & _T_269;
  assign _T_271 = _T_255 | _T_270;
  assign _T_272 = _T_242[0];
  assign _T_273 = io_out_1_a_bits_address[0];
  assign _T_275 = _T_273 == 1'h0;
  assign _T_276 = _T_260 & _T_275;
  assign _T_277 = _T_272 & _T_276;
  assign _T_278 = _T_262 | _T_277;
  assign _T_279 = _T_260 & _T_273;
  assign _T_280 = _T_272 & _T_279;
  assign _T_281 = _T_262 | _T_280;
  assign _T_282 = _T_263 & _T_275;
  assign _T_283 = _T_272 & _T_282;
  assign _T_284 = _T_265 | _T_283;
  assign _T_285 = _T_263 & _T_273;
  assign _T_286 = _T_272 & _T_285;
  assign _T_287 = _T_265 | _T_286;
  assign _T_288 = _T_266 & _T_275;
  assign _T_289 = _T_272 & _T_288;
  assign _T_290 = _T_268 | _T_289;
  assign _T_291 = _T_266 & _T_273;
  assign _T_292 = _T_272 & _T_291;
  assign _T_293 = _T_268 | _T_292;
  assign _T_294 = _T_269 & _T_275;
  assign _T_295 = _T_272 & _T_294;
  assign _T_296 = _T_271 | _T_295;
  assign _T_297 = _T_269 & _T_273;
  assign _T_298 = _T_272 & _T_297;
  assign _T_299 = _T_271 | _T_298;
  assign _T_300 = {_T_281,_T_278};
  assign _T_301 = {_T_287,_T_284};
  assign _T_302 = {_T_301,_T_300};
  assign _T_303 = {_T_293,_T_290};
  assign _T_304 = {_T_299,_T_296};
  assign _T_305 = {_T_304,_T_303};
  assign _T_306 = {_T_305,_T_302};
  assign _T_313 = _T_207 ? io_in_1_a_bits_mask : _T_309_0;
  assign _GEN_6 = _T_235 ? _T_313 : _T_309_0;
  assign _T_319 = {io_in_1_a_bits_mask,_T_313};
  assign _T_322 = _T_185 ? _T_319 : 8'hff;
  assign _T_323 = _T_306 & _T_322;
  assign Repeater_clock = clock;
  assign Repeater_reset = reset;
  assign Repeater_io_repeat = _T_405;
  assign Repeater_io_enq_valid = io_out_1_d_valid;
  assign Repeater_io_enq_bits_opcode = io_out_1_d_bits_opcode;
  assign Repeater_io_enq_bits_param = io_out_1_d_bits_param;
  assign Repeater_io_enq_bits_size = io_out_1_d_bits_size;
  assign Repeater_io_enq_bits_source = io_out_1_d_bits_source;
  assign Repeater_io_enq_bits_sink = io_out_1_d_bits_sink;
  assign Repeater_io_enq_bits_data = io_out_1_d_bits_data;
  assign Repeater_io_enq_bits_error = io_out_1_d_bits_error;
  assign Repeater_io_deq_ready = io_in_1_d_ready;
  assign _T_326_valid = Repeater_io_deq_valid;
  assign _T_326_bits_opcode = Repeater_io_deq_bits_opcode;
  assign _T_326_bits_param = Repeater_io_deq_bits_param;
  assign _T_326_bits_size = Repeater_io_deq_bits_size;
  assign _T_326_bits_source = Repeater_io_deq_bits_source;
  assign _T_326_bits_sink = Repeater_io_deq_bits_sink;
  assign _T_326_bits_error = Repeater_io_deq_bits_error;
  assign _T_330 = Repeater_io_deq_bits_data[63:32];
  assign _T_331 = io_out_1_d_bits_data[31:0];
  assign _T_332 = {_T_330,_T_331};
  assign _T_333 = _T_326_bits_opcode[0];
  assign _T_336 = 18'h7 << _T_326_bits_size;
  assign _T_337 = _T_336[2:0];
  assign _T_338 = ~ _T_337;
  assign _T_339 = _T_338[2:2];
  assign _T_344 = _T_342 == 1'h0;
  assign _T_345 = _T_342 == _T_339;
  assign _T_347 = _T_333 == 1'h0;
  assign _T_348 = _T_345 | _T_347;
  assign _T_349 = io_in_1_d_ready & io_in_1_d_valid;
  assign _T_351 = _T_342 + 1'h1;
  assign _T_352 = _T_351[0:0];
  assign _GEN_7 = _T_348 ? 1'h0 : _T_352;
  assign _GEN_8 = _T_349 ? _GEN_7 : _T_342;
  assign _T_378 = io_in_1_a_bits_address[2];
  assign _GEN_9 = 5'h0 == io_in_1_a_bits_source ? _T_378 : _T_357_0;
  assign _GEN_10 = 5'h1 == io_in_1_a_bits_source ? _T_378 : _T_357_1;
  assign _GEN_11 = 5'h2 == io_in_1_a_bits_source ? _T_378 : _T_357_2;
  assign _GEN_12 = 5'h3 == io_in_1_a_bits_source ? _T_378 : _T_357_3;
  assign _GEN_13 = 5'h4 == io_in_1_a_bits_source ? _T_378 : _T_357_4;
  assign _GEN_14 = 5'h5 == io_in_1_a_bits_source ? _T_378 : _T_357_5;
  assign _GEN_15 = 5'h6 == io_in_1_a_bits_source ? _T_378 : _T_357_6;
  assign _GEN_16 = 5'h7 == io_in_1_a_bits_source ? _T_378 : _T_357_7;
  assign _GEN_17 = 5'h8 == io_in_1_a_bits_source ? _T_378 : _T_357_8;
  assign _GEN_18 = 5'h9 == io_in_1_a_bits_source ? _T_378 : _T_357_9;
  assign _GEN_19 = 5'ha == io_in_1_a_bits_source ? _T_378 : _T_357_10;
  assign _GEN_20 = 5'hb == io_in_1_a_bits_source ? _T_378 : _T_357_11;
  assign _GEN_21 = 5'hc == io_in_1_a_bits_source ? _T_378 : _T_357_12;
  assign _GEN_22 = 5'hd == io_in_1_a_bits_source ? _T_378 : _T_357_13;
  assign _GEN_23 = 5'he == io_in_1_a_bits_source ? _T_378 : _T_357_14;
  assign _GEN_24 = 5'hf == io_in_1_a_bits_source ? _T_378 : _T_357_15;
  assign _GEN_25 = 5'h10 == io_in_1_a_bits_source ? _T_378 : _T_357_16;
  assign _GEN_26 = 5'h11 == io_in_1_a_bits_source ? _T_378 : _T_357_17;
  assign _GEN_27 = _T_215 ? _GEN_9 : _T_357_0;
  assign _GEN_28 = _T_215 ? _GEN_10 : _T_357_1;
  assign _GEN_29 = _T_215 ? _GEN_11 : _T_357_2;
  assign _GEN_30 = _T_215 ? _GEN_12 : _T_357_3;
  assign _GEN_31 = _T_215 ? _GEN_13 : _T_357_4;
  assign _GEN_32 = _T_215 ? _GEN_14 : _T_357_5;
  assign _GEN_33 = _T_215 ? _GEN_15 : _T_357_6;
  assign _GEN_34 = _T_215 ? _GEN_16 : _T_357_7;
  assign _GEN_35 = _T_215 ? _GEN_17 : _T_357_8;
  assign _GEN_36 = _T_215 ? _GEN_18 : _T_357_9;
  assign _GEN_37 = _T_215 ? _GEN_19 : _T_357_10;
  assign _GEN_38 = _T_215 ? _GEN_20 : _T_357_11;
  assign _GEN_39 = _T_215 ? _GEN_21 : _T_357_12;
  assign _GEN_40 = _T_215 ? _GEN_22 : _T_357_13;
  assign _GEN_41 = _T_215 ? _GEN_23 : _T_357_14;
  assign _GEN_42 = _T_215 ? _GEN_24 : _T_357_15;
  assign _GEN_43 = _T_215 ? _GEN_25 : _T_357_16;
  assign _GEN_44 = _T_215 ? _GEN_26 : _T_357_17;
  assign _GEN_45 = 5'h1 == _T_326_bits_source ? _T_357_1 : _T_357_0;
  assign _GEN_46 = 5'h2 == _T_326_bits_source ? _T_357_2 : _GEN_45;
  assign _GEN_47 = 5'h3 == _T_326_bits_source ? _T_357_3 : _GEN_46;
  assign _GEN_48 = 5'h4 == _T_326_bits_source ? _T_357_4 : _GEN_47;
  assign _GEN_49 = 5'h5 == _T_326_bits_source ? _T_357_5 : _GEN_48;
  assign _GEN_50 = 5'h6 == _T_326_bits_source ? _T_357_6 : _GEN_49;
  assign _GEN_51 = 5'h7 == _T_326_bits_source ? _T_357_7 : _GEN_50;
  assign _GEN_52 = 5'h8 == _T_326_bits_source ? _T_357_8 : _GEN_51;
  assign _GEN_53 = 5'h9 == _T_326_bits_source ? _T_357_9 : _GEN_52;
  assign _GEN_54 = 5'ha == _T_326_bits_source ? _T_357_10 : _GEN_53;
  assign _GEN_55 = 5'hb == _T_326_bits_source ? _T_357_11 : _GEN_54;
  assign _GEN_56 = 5'hc == _T_326_bits_source ? _T_357_12 : _GEN_55;
  assign _GEN_57 = 5'hd == _T_326_bits_source ? _T_357_13 : _GEN_56;
  assign _GEN_58 = 5'he == _T_326_bits_source ? _T_357_14 : _GEN_57;
  assign _GEN_59 = 5'hf == _T_326_bits_source ? _T_357_15 : _GEN_58;
  assign _GEN_60 = 5'h10 == _T_326_bits_source ? _T_357_16 : _GEN_59;
  assign _GEN_61 = 5'h11 == _T_326_bits_source ? _T_357_17 : _GEN_60;
  assign _GEN_62 = _T_344 ? _GEN_61 : _T_389;
  assign _T_391 = ~ _T_339;
  assign _T_392 = _GEN_62 & _T_391;
  assign _T_393 = _T_392 | _T_342;
  assign _T_394 = _T_332[31:0];
  assign _T_395 = _T_332[63:32];
  assign _GEN_63 = _T_393 ? _T_395 : _T_394;
  assign _T_405 = _T_348 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_194 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_226_0 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_309_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_342 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_357_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_357_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_357_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_357_3 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_357_4 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_357_5 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_357_6 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_357_7 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_357_8 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_357_9 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_357_10 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_357_11 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_357_12 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_357_13 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_357_14 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_357_15 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_357_16 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_357_17 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_389 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_194 <= 1'h0;
    end else begin
      if (_T_215) begin
        if (_T_200) begin
          _T_194 <= 1'h0;
        end else begin
          _T_194 <= _T_218;
        end
      end
    end
    if (_T_235) begin
      if (_T_207) begin
        _T_226_0 <= io_in_1_a_bits_data;
      end
    end
    if (_T_235) begin
      if (_T_207) begin
        _T_309_0 <= io_in_1_a_bits_mask;
      end
    end
    if (reset) begin
      _T_342 <= 1'h0;
    end else begin
      if (_T_349) begin
        if (_T_348) begin
          _T_342 <= 1'h0;
        end else begin
          _T_342 <= _T_352;
        end
      end
    end
    if (_T_215) begin
      if (5'h0 == io_in_1_a_bits_source) begin
        _T_357_0 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h1 == io_in_1_a_bits_source) begin
        _T_357_1 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h2 == io_in_1_a_bits_source) begin
        _T_357_2 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h3 == io_in_1_a_bits_source) begin
        _T_357_3 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h4 == io_in_1_a_bits_source) begin
        _T_357_4 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h5 == io_in_1_a_bits_source) begin
        _T_357_5 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h6 == io_in_1_a_bits_source) begin
        _T_357_6 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h7 == io_in_1_a_bits_source) begin
        _T_357_7 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h8 == io_in_1_a_bits_source) begin
        _T_357_8 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h9 == io_in_1_a_bits_source) begin
        _T_357_9 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'ha == io_in_1_a_bits_source) begin
        _T_357_10 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'hb == io_in_1_a_bits_source) begin
        _T_357_11 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'hc == io_in_1_a_bits_source) begin
        _T_357_12 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'hd == io_in_1_a_bits_source) begin
        _T_357_13 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'he == io_in_1_a_bits_source) begin
        _T_357_14 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'hf == io_in_1_a_bits_source) begin
        _T_357_15 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h10 == io_in_1_a_bits_source) begin
        _T_357_16 <= _T_378;
      end
    end
    if (_T_215) begin
      if (5'h11 == io_in_1_a_bits_source) begin
        _T_357_17 <= _T_378;
      end
    end
    if (_T_344) begin
      if (5'h11 == _T_326_bits_source) begin
        _T_389 <= _T_357_17;
      end else begin
        if (5'h10 == _T_326_bits_source) begin
          _T_389 <= _T_357_16;
        end else begin
          if (5'hf == _T_326_bits_source) begin
            _T_389 <= _T_357_15;
          end else begin
            if (5'he == _T_326_bits_source) begin
              _T_389 <= _T_357_14;
            end else begin
              if (5'hd == _T_326_bits_source) begin
                _T_389 <= _T_357_13;
              end else begin
                if (5'hc == _T_326_bits_source) begin
                  _T_389 <= _T_357_12;
                end else begin
                  if (5'hb == _T_326_bits_source) begin
                    _T_389 <= _T_357_11;
                  end else begin
                    if (5'ha == _T_326_bits_source) begin
                      _T_389 <= _T_357_10;
                    end else begin
                      if (5'h9 == _T_326_bits_source) begin
                        _T_389 <= _T_357_9;
                      end else begin
                        if (5'h8 == _T_326_bits_source) begin
                          _T_389 <= _T_357_8;
                        end else begin
                          if (5'h7 == _T_326_bits_source) begin
                            _T_389 <= _T_357_7;
                          end else begin
                            if (5'h6 == _T_326_bits_source) begin
                              _T_389 <= _T_357_6;
                            end else begin
                              if (5'h5 == _T_326_bits_source) begin
                                _T_389 <= _T_357_5;
                              end else begin
                                if (5'h4 == _T_326_bits_source) begin
                                  _T_389 <= _T_357_4;
                                end else begin
                                  if (5'h3 == _T_326_bits_source) begin
                                    _T_389 <= _T_357_3;
                                  end else begin
                                    if (5'h2 == _T_326_bits_source) begin
                                      _T_389 <= _T_357_2;
                                    end else begin
                                      if (5'h1 == _T_326_bits_source) begin
                                        _T_389 <= _T_357_1;
                                      end else begin
                                        _T_389 <= _T_357_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module TLSplitter(
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [2:0]  io_in_1_a_bits_param,
  input  [3:0]  io_in_1_a_bits_size,
  input  [3:0]  io_in_1_a_bits_source,
  input  [31:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [3:0]  io_in_1_d_bits_size,
  output [3:0]  io_in_1_d_bits_source,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input         io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output        io_in_0_d_bits_source,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [2:0]  io_out_1_a_bits_param,
  output [3:0]  io_out_1_a_bits_size,
  output [3:0]  io_out_1_a_bits_source,
  output [31:0] io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [3:0]  io_out_1_d_bits_size,
  input  [3:0]  io_out_1_d_bits_source,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input         io_out_0_d_bits_source,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  assign io_in_1_a_ready = io_out_1_a_ready;
  assign io_in_1_d_valid = io_out_1_d_valid;
  assign io_in_1_d_bits_opcode = io_out_1_d_bits_opcode;
  assign io_in_1_d_bits_size = io_out_1_d_bits_size;
  assign io_in_1_d_bits_source = io_out_1_d_bits_source;
  assign io_in_0_a_ready = io_out_0_a_ready;
  assign io_in_0_d_valid = io_out_0_d_valid;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_d_bits_error = io_out_0_d_bits_error;
  assign io_out_1_a_valid = io_in_1_a_valid;
  assign io_out_1_a_bits_opcode = io_in_1_a_bits_opcode;
  assign io_out_1_a_bits_param = io_in_1_a_bits_param;
  assign io_out_1_a_bits_size = io_in_1_a_bits_size;
  assign io_out_1_a_bits_source = io_in_1_a_bits_source;
  assign io_out_1_a_bits_address = io_in_1_a_bits_address;
  assign io_out_1_a_bits_mask = io_in_1_a_bits_mask;
  assign io_out_1_a_bits_data = io_in_1_a_bits_data;
  assign io_out_1_d_ready = io_in_1_d_ready;
  assign io_out_0_a_valid = io_in_0_a_valid;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_param = io_in_0_a_bits_param;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address;
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = io_in_0_d_ready;
endmodule
module TLFIFOFixer(
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input         io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output        io_in_0_d_bits_source,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input         io_out_0_d_bits_source,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  assign io_in_0_a_ready = io_out_0_a_ready;
  assign io_in_0_d_valid = io_out_0_d_valid;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_d_bits_error = io_out_0_d_bits_error;
  assign io_out_0_a_valid = io_in_0_a_valid;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_param = io_in_0_a_bits_param;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address;
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = io_in_0_d_ready;
endmodule
module TLFIFOFixer_1(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input  [3:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output [3:0]  io_in_0_d_bits_source,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output [3:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input  [3:0]  io_out_0_d_bits_source
);
  wire [32:0] _T_92;
  wire [32:0] _T_103;
  wire [32:0] _T_104;
  wire  _T_106;
  wire [31:0] _T_109;
  wire [32:0] _T_110;
  wire [32:0] _T_112;
  wire [32:0] _T_113;
  wire  _T_115;
  wire [31:0] _T_118;
  wire [32:0] _T_119;
  wire [32:0] _T_121;
  wire [32:0] _T_122;
  wire  _T_124;
  wire [31:0] _T_127;
  wire [32:0] _T_128;
  wire [32:0] _T_130;
  wire [32:0] _T_131;
  wire  _T_133;
  wire [31:0] _T_136;
  wire [32:0] _T_137;
  wire [32:0] _T_139;
  wire [32:0] _T_140;
  wire  _T_142;
  wire [31:0] _T_145;
  wire [32:0] _T_146;
  wire [32:0] _T_148;
  wire [32:0] _T_149;
  wire  _T_151;
  wire [31:0] _T_154;
  wire [32:0] _T_155;
  wire [32:0] _T_157;
  wire [32:0] _T_158;
  wire  _T_160;
  wire [1:0] _T_166;
  wire [2:0] _T_168;
  wire [1:0] _T_170;
  wire [2:0] _T_172;
  wire [2:0] _T_174;
  wire [2:0] _T_176;
  wire [1:0] _GEN_70;
  wire [1:0] _T_177;
  wire [2:0] _GEN_71;
  wire [2:0] _T_178;
  wire [2:0] _GEN_72;
  wire [2:0] _T_179;
  wire [2:0] _T_180;
  wire [2:0] _T_181;
  wire [2:0] _T_182;
  wire  _T_186;
  wire  _T_187;
  wire [26:0] _T_190;
  wire [11:0] _T_191;
  wire [11:0] _T_192;
  wire [9:0] _T_193;
  wire  _T_194;
  wire  _T_196;
  wire [9:0] _T_198;
  reg [9:0] _T_201;
  reg [31:0] _RAND_0;
  wire [10:0] _T_203;
  wire [10:0] _T_204;
  wire [9:0] _T_205;
  wire  _T_207;
  wire [9:0] _T_216;
  wire [9:0] _GEN_2;
  wire  _T_217;
  wire [26:0] _T_220;
  wire [11:0] _T_221;
  wire [11:0] _T_222;
  wire [9:0] _T_223;
  wire  _T_224;
  wire [9:0] _T_226;
  reg [9:0] _T_229;
  reg [31:0] _RAND_1;
  wire [10:0] _T_231;
  wire [10:0] _T_232;
  wire [9:0] _T_233;
  wire  _T_235;
  wire [9:0] _T_244;
  wire [9:0] _GEN_3;
  wire  _T_246;
  wire  _T_247;
  reg  _T_321_0;
  reg [31:0] _RAND_2;
  reg  _T_321_1;
  reg [31:0] _RAND_3;
  reg  _T_321_2;
  reg [31:0] _RAND_4;
  reg  _T_321_3;
  reg [31:0] _RAND_5;
  reg  _T_321_4;
  reg [31:0] _RAND_6;
  reg  _T_321_5;
  reg [31:0] _RAND_7;
  reg  _T_321_6;
  reg [31:0] _RAND_8;
  reg  _T_321_7;
  reg [31:0] _RAND_9;
  reg  _T_321_8;
  reg [31:0] _RAND_10;
  reg  _T_321_9;
  reg [31:0] _RAND_11;
  reg  _T_321_10;
  reg [31:0] _RAND_12;
  reg  _T_321_11;
  reg [31:0] _RAND_13;
  reg  _T_321_12;
  reg [31:0] _RAND_14;
  reg  _T_321_13;
  reg [31:0] _RAND_15;
  reg  _T_321_14;
  reg [31:0] _RAND_16;
  reg  _T_321_15;
  reg [31:0] _RAND_17;
  wire  _T_375;
  wire  _GEN_4;
  wire  _GEN_5;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _T_381;
  wire  _T_382;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _T_390;
  wire  _T_392;
  wire  _T_400;
  reg [2:0] _T_405;
  reg [31:0] _RAND_18;
  wire [2:0] _GEN_68;
  wire  _T_406;
  wire  _T_407;
  wire  _T_408;
  wire  _T_409;
  wire  _T_410;
  wire  _T_411;
  wire  _T_412;
  wire  _T_413;
  wire  _T_414;
  wire  _T_415;
  wire  _T_416;
  wire  _T_417;
  wire  _T_431;
  reg [2:0] _T_436;
  reg [31:0] _RAND_19;
  wire [2:0] _GEN_69;
  wire  _T_437;
  wire  _T_438;
  wire  _T_439;
  wire  _T_440;
  wire  _T_441;
  wire  _T_442;
  wire  _T_443;
  wire  _T_444;
  wire  _T_445;
  wire  _T_446;
  wire  _T_447;
  wire  _T_448;
  wire  _T_451;
  wire  _T_453;
  wire  _T_455;
  wire  _T_459;
  assign io_in_0_a_ready = _T_459;
  assign io_in_0_d_valid = io_out_0_d_valid;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_out_0_a_valid = _T_455;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_param = io_in_0_a_bits_param;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address;
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = io_in_0_d_ready;
  assign _T_92 = {1'b0,$signed(io_in_0_a_bits_address)};
  assign _T_103 = $signed(_T_92) & $signed(33'sha6011000);
  assign _T_104 = $signed(_T_103);
  assign _T_106 = $signed(_T_104) == $signed(33'sh0);
  assign _T_109 = io_in_0_a_bits_address ^ 32'h4000000;
  assign _T_110 = {1'b0,$signed(_T_109)};
  assign _T_112 = $signed(_T_110) & $signed(33'sha4000000);
  assign _T_113 = $signed(_T_112);
  assign _T_115 = $signed(_T_113) == $signed(33'sh0);
  assign _T_118 = io_in_0_a_bits_address ^ 32'h10000;
  assign _T_119 = {1'b0,$signed(_T_118)};
  assign _T_121 = $signed(_T_119) & $signed(33'sha6010000);
  assign _T_122 = $signed(_T_121);
  assign _T_124 = $signed(_T_122) == $signed(33'sh0);
  assign _T_127 = io_in_0_a_bits_address ^ 32'h20000000;
  assign _T_128 = {1'b0,$signed(_T_127)};
  assign _T_130 = $signed(_T_128) & $signed(33'sha0000000);
  assign _T_131 = $signed(_T_130);
  assign _T_133 = $signed(_T_131) == $signed(33'sh0);
  assign _T_136 = io_in_0_a_bits_address ^ 32'h80000000;
  assign _T_137 = {1'b0,$signed(_T_136)};
  assign _T_139 = $signed(_T_137) & $signed(33'sha6010000);
  assign _T_140 = $signed(_T_139);
  assign _T_142 = $signed(_T_140) == $signed(33'sh0);
  assign _T_145 = io_in_0_a_bits_address ^ 32'h2000000;
  assign _T_146 = {1'b0,$signed(_T_145)};
  assign _T_148 = $signed(_T_146) & $signed(33'sha6010000);
  assign _T_149 = $signed(_T_148);
  assign _T_151 = $signed(_T_149) == $signed(33'sh0);
  assign _T_154 = io_in_0_a_bits_address ^ 32'h1000;
  assign _T_155 = {1'b0,$signed(_T_154)};
  assign _T_157 = $signed(_T_155) & $signed(33'sha6011000);
  assign _T_158 = $signed(_T_157);
  assign _T_160 = $signed(_T_158) == $signed(33'sh0);
  assign _T_166 = _T_133 ? 2'h2 : 2'h0;
  assign _T_168 = _T_106 ? 3'h5 : 3'h0;
  assign _T_170 = _T_151 ? 2'h3 : 2'h0;
  assign _T_172 = _T_142 ? 3'h7 : 3'h0;
  assign _T_174 = _T_124 ? 3'h6 : 3'h0;
  assign _T_176 = _T_160 ? 3'h4 : 3'h0;
  assign _GEN_70 = {{1'd0}, _T_115};
  assign _T_177 = _GEN_70 | _T_166;
  assign _GEN_71 = {{1'd0}, _T_177};
  assign _T_178 = _GEN_71 | _T_168;
  assign _GEN_72 = {{1'd0}, _T_170};
  assign _T_179 = _T_178 | _GEN_72;
  assign _T_180 = _T_179 | _T_172;
  assign _T_181 = _T_180 | _T_174;
  assign _T_182 = _T_181 | _T_176;
  assign _T_186 = _T_182 == 3'h0;
  assign _T_187 = io_in_0_a_ready & io_in_0_a_valid;
  assign _T_190 = 27'hfff << io_in_0_a_bits_size;
  assign _T_191 = _T_190[11:0];
  assign _T_192 = ~ _T_191;
  assign _T_193 = _T_192[11:2];
  assign _T_194 = io_in_0_a_bits_opcode[2];
  assign _T_196 = _T_194 == 1'h0;
  assign _T_198 = _T_196 ? _T_193 : 10'h0;
  assign _T_203 = _T_201 - 10'h1;
  assign _T_204 = $unsigned(_T_203);
  assign _T_205 = _T_204[9:0];
  assign _T_207 = _T_201 == 10'h0;
  assign _T_216 = _T_207 ? _T_198 : _T_205;
  assign _GEN_2 = _T_187 ? _T_216 : _T_201;
  assign _T_217 = io_out_0_d_ready & io_out_0_d_valid;
  assign _T_220 = 27'hfff << io_out_0_d_bits_size;
  assign _T_221 = _T_220[11:0];
  assign _T_222 = ~ _T_221;
  assign _T_223 = _T_222[11:2];
  assign _T_224 = io_out_0_d_bits_opcode[0];
  assign _T_226 = _T_224 ? _T_223 : 10'h0;
  assign _T_231 = _T_229 - 10'h1;
  assign _T_232 = $unsigned(_T_231);
  assign _T_233 = _T_232[9:0];
  assign _T_235 = _T_229 == 10'h0;
  assign _T_244 = _T_235 ? _T_226 : _T_233;
  assign _GEN_3 = _T_217 ? _T_244 : _T_229;
  assign _T_246 = io_out_0_d_bits_opcode != 3'h6;
  assign _T_247 = _T_235 & _T_246;
  assign _T_375 = _T_207 & _T_187;
  assign _GEN_4 = 4'h0 == io_in_0_a_bits_source ? 1'h1 : _T_321_0;
  assign _GEN_5 = 4'h1 == io_in_0_a_bits_source ? 1'h1 : _T_321_1;
  assign _GEN_6 = 4'h2 == io_in_0_a_bits_source ? 1'h1 : _T_321_2;
  assign _GEN_7 = 4'h3 == io_in_0_a_bits_source ? 1'h1 : _T_321_3;
  assign _GEN_8 = 4'h4 == io_in_0_a_bits_source ? 1'h1 : _T_321_4;
  assign _GEN_9 = 4'h5 == io_in_0_a_bits_source ? 1'h1 : _T_321_5;
  assign _GEN_10 = 4'h6 == io_in_0_a_bits_source ? 1'h1 : _T_321_6;
  assign _GEN_11 = 4'h7 == io_in_0_a_bits_source ? 1'h1 : _T_321_7;
  assign _GEN_12 = 4'h8 == io_in_0_a_bits_source ? 1'h1 : _T_321_8;
  assign _GEN_13 = 4'h9 == io_in_0_a_bits_source ? 1'h1 : _T_321_9;
  assign _GEN_14 = 4'ha == io_in_0_a_bits_source ? 1'h1 : _T_321_10;
  assign _GEN_15 = 4'hb == io_in_0_a_bits_source ? 1'h1 : _T_321_11;
  assign _GEN_16 = 4'hc == io_in_0_a_bits_source ? 1'h1 : _T_321_12;
  assign _GEN_17 = 4'hd == io_in_0_a_bits_source ? 1'h1 : _T_321_13;
  assign _GEN_18 = 4'he == io_in_0_a_bits_source ? 1'h1 : _T_321_14;
  assign _GEN_19 = 4'hf == io_in_0_a_bits_source ? 1'h1 : _T_321_15;
  assign _GEN_20 = _T_375 ? _GEN_4 : _T_321_0;
  assign _GEN_21 = _T_375 ? _GEN_5 : _T_321_1;
  assign _GEN_22 = _T_375 ? _GEN_6 : _T_321_2;
  assign _GEN_23 = _T_375 ? _GEN_7 : _T_321_3;
  assign _GEN_24 = _T_375 ? _GEN_8 : _T_321_4;
  assign _GEN_25 = _T_375 ? _GEN_9 : _T_321_5;
  assign _GEN_26 = _T_375 ? _GEN_10 : _T_321_6;
  assign _GEN_27 = _T_375 ? _GEN_11 : _T_321_7;
  assign _GEN_28 = _T_375 ? _GEN_12 : _T_321_8;
  assign _GEN_29 = _T_375 ? _GEN_13 : _T_321_9;
  assign _GEN_30 = _T_375 ? _GEN_14 : _T_321_10;
  assign _GEN_31 = _T_375 ? _GEN_15 : _T_321_11;
  assign _GEN_32 = _T_375 ? _GEN_16 : _T_321_12;
  assign _GEN_33 = _T_375 ? _GEN_17 : _T_321_13;
  assign _GEN_34 = _T_375 ? _GEN_18 : _T_321_14;
  assign _GEN_35 = _T_375 ? _GEN_19 : _T_321_15;
  assign _T_381 = io_in_0_d_ready & io_in_0_d_valid;
  assign _T_382 = _T_247 & _T_381;
  assign _GEN_36 = 4'h0 == io_in_0_d_bits_source ? 1'h0 : _GEN_20;
  assign _GEN_37 = 4'h1 == io_in_0_d_bits_source ? 1'h0 : _GEN_21;
  assign _GEN_38 = 4'h2 == io_in_0_d_bits_source ? 1'h0 : _GEN_22;
  assign _GEN_39 = 4'h3 == io_in_0_d_bits_source ? 1'h0 : _GEN_23;
  assign _GEN_40 = 4'h4 == io_in_0_d_bits_source ? 1'h0 : _GEN_24;
  assign _GEN_41 = 4'h5 == io_in_0_d_bits_source ? 1'h0 : _GEN_25;
  assign _GEN_42 = 4'h6 == io_in_0_d_bits_source ? 1'h0 : _GEN_26;
  assign _GEN_43 = 4'h7 == io_in_0_d_bits_source ? 1'h0 : _GEN_27;
  assign _GEN_44 = 4'h8 == io_in_0_d_bits_source ? 1'h0 : _GEN_28;
  assign _GEN_45 = 4'h9 == io_in_0_d_bits_source ? 1'h0 : _GEN_29;
  assign _GEN_46 = 4'ha == io_in_0_d_bits_source ? 1'h0 : _GEN_30;
  assign _GEN_47 = 4'hb == io_in_0_d_bits_source ? 1'h0 : _GEN_31;
  assign _GEN_48 = 4'hc == io_in_0_d_bits_source ? 1'h0 : _GEN_32;
  assign _GEN_49 = 4'hd == io_in_0_d_bits_source ? 1'h0 : _GEN_33;
  assign _GEN_50 = 4'he == io_in_0_d_bits_source ? 1'h0 : _GEN_34;
  assign _GEN_51 = 4'hf == io_in_0_d_bits_source ? 1'h0 : _GEN_35;
  assign _GEN_52 = _T_382 ? _GEN_36 : _GEN_20;
  assign _GEN_53 = _T_382 ? _GEN_37 : _GEN_21;
  assign _GEN_54 = _T_382 ? _GEN_38 : _GEN_22;
  assign _GEN_55 = _T_382 ? _GEN_39 : _GEN_23;
  assign _GEN_56 = _T_382 ? _GEN_40 : _GEN_24;
  assign _GEN_57 = _T_382 ? _GEN_41 : _GEN_25;
  assign _GEN_58 = _T_382 ? _GEN_42 : _GEN_26;
  assign _GEN_59 = _T_382 ? _GEN_43 : _GEN_27;
  assign _GEN_60 = _T_382 ? _GEN_44 : _GEN_28;
  assign _GEN_61 = _T_382 ? _GEN_45 : _GEN_29;
  assign _GEN_62 = _T_382 ? _GEN_46 : _GEN_30;
  assign _GEN_63 = _T_382 ? _GEN_47 : _GEN_31;
  assign _GEN_64 = _T_382 ? _GEN_48 : _GEN_32;
  assign _GEN_65 = _T_382 ? _GEN_49 : _GEN_33;
  assign _GEN_66 = _T_382 ? _GEN_50 : _GEN_34;
  assign _GEN_67 = _T_382 ? _GEN_51 : _GEN_35;
  assign _T_390 = io_in_0_a_bits_source[3:3];
  assign _T_392 = _T_390 == 1'h0;
  assign _T_400 = _T_187 & _T_392;
  assign _GEN_68 = _T_400 ? _T_182 : _T_405;
  assign _T_406 = _T_392 & _T_207;
  assign _T_407 = _T_321_0 | _T_321_1;
  assign _T_408 = _T_407 | _T_321_2;
  assign _T_409 = _T_408 | _T_321_3;
  assign _T_410 = _T_409 | _T_321_4;
  assign _T_411 = _T_410 | _T_321_5;
  assign _T_412 = _T_411 | _T_321_6;
  assign _T_413 = _T_412 | _T_321_7;
  assign _T_414 = _T_406 & _T_413;
  assign _T_415 = _T_405 != _T_182;
  assign _T_416 = _T_186 | _T_415;
  assign _T_417 = _T_414 & _T_416;
  assign _T_431 = _T_187 & _T_390;
  assign _GEN_69 = _T_431 ? _T_182 : _T_436;
  assign _T_437 = _T_390 & _T_207;
  assign _T_438 = _T_321_8 | _T_321_9;
  assign _T_439 = _T_438 | _T_321_10;
  assign _T_440 = _T_439 | _T_321_11;
  assign _T_441 = _T_440 | _T_321_12;
  assign _T_442 = _T_441 | _T_321_13;
  assign _T_443 = _T_442 | _T_321_14;
  assign _T_444 = _T_443 | _T_321_15;
  assign _T_445 = _T_437 & _T_444;
  assign _T_446 = _T_436 != _T_182;
  assign _T_447 = _T_186 | _T_446;
  assign _T_448 = _T_445 & _T_447;
  assign _T_451 = _T_417 | _T_448;
  assign _T_453 = _T_451 == 1'h0;
  assign _T_455 = io_in_0_a_valid & _T_453;
  assign _T_459 = io_out_0_a_ready & _T_453;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_201 = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_229 = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_321_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_321_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_321_2 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_321_3 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_321_4 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_321_5 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_321_6 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_321_7 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_321_8 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_321_9 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_321_10 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_321_11 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_321_12 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_321_13 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_321_14 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_321_15 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_405 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_436 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_201 <= 10'h0;
    end else begin
      if (_T_187) begin
        if (_T_207) begin
          if (_T_196) begin
            _T_201 <= _T_193;
          end else begin
            _T_201 <= 10'h0;
          end
        end else begin
          _T_201 <= _T_205;
        end
      end
    end
    if (reset) begin
      _T_229 <= 10'h0;
    end else begin
      if (_T_217) begin
        if (_T_235) begin
          if (_T_224) begin
            _T_229 <= _T_223;
          end else begin
            _T_229 <= 10'h0;
          end
        end else begin
          _T_229 <= _T_233;
        end
      end
    end
    if (reset) begin
      _T_321_0 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h0 == io_in_0_d_bits_source) begin
          _T_321_0 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h0 == io_in_0_a_bits_source) begin
              _T_321_0 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h0 == io_in_0_a_bits_source) begin
            _T_321_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_1 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h1 == io_in_0_d_bits_source) begin
          _T_321_1 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h1 == io_in_0_a_bits_source) begin
              _T_321_1 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h1 == io_in_0_a_bits_source) begin
            _T_321_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_2 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h2 == io_in_0_d_bits_source) begin
          _T_321_2 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h2 == io_in_0_a_bits_source) begin
              _T_321_2 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h2 == io_in_0_a_bits_source) begin
            _T_321_2 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_3 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h3 == io_in_0_d_bits_source) begin
          _T_321_3 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h3 == io_in_0_a_bits_source) begin
              _T_321_3 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h3 == io_in_0_a_bits_source) begin
            _T_321_3 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_4 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h4 == io_in_0_d_bits_source) begin
          _T_321_4 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h4 == io_in_0_a_bits_source) begin
              _T_321_4 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h4 == io_in_0_a_bits_source) begin
            _T_321_4 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_5 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h5 == io_in_0_d_bits_source) begin
          _T_321_5 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h5 == io_in_0_a_bits_source) begin
              _T_321_5 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h5 == io_in_0_a_bits_source) begin
            _T_321_5 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_6 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h6 == io_in_0_d_bits_source) begin
          _T_321_6 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h6 == io_in_0_a_bits_source) begin
              _T_321_6 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h6 == io_in_0_a_bits_source) begin
            _T_321_6 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_7 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h7 == io_in_0_d_bits_source) begin
          _T_321_7 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h7 == io_in_0_a_bits_source) begin
              _T_321_7 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h7 == io_in_0_a_bits_source) begin
            _T_321_7 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_8 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h8 == io_in_0_d_bits_source) begin
          _T_321_8 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h8 == io_in_0_a_bits_source) begin
              _T_321_8 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h8 == io_in_0_a_bits_source) begin
            _T_321_8 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_9 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'h9 == io_in_0_d_bits_source) begin
          _T_321_9 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'h9 == io_in_0_a_bits_source) begin
              _T_321_9 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'h9 == io_in_0_a_bits_source) begin
            _T_321_9 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_10 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'ha == io_in_0_d_bits_source) begin
          _T_321_10 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'ha == io_in_0_a_bits_source) begin
              _T_321_10 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'ha == io_in_0_a_bits_source) begin
            _T_321_10 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_11 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'hb == io_in_0_d_bits_source) begin
          _T_321_11 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'hb == io_in_0_a_bits_source) begin
              _T_321_11 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'hb == io_in_0_a_bits_source) begin
            _T_321_11 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_12 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'hc == io_in_0_d_bits_source) begin
          _T_321_12 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'hc == io_in_0_a_bits_source) begin
              _T_321_12 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'hc == io_in_0_a_bits_source) begin
            _T_321_12 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_13 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'hd == io_in_0_d_bits_source) begin
          _T_321_13 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'hd == io_in_0_a_bits_source) begin
              _T_321_13 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'hd == io_in_0_a_bits_source) begin
            _T_321_13 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_14 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'he == io_in_0_d_bits_source) begin
          _T_321_14 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'he == io_in_0_a_bits_source) begin
              _T_321_14 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'he == io_in_0_a_bits_source) begin
            _T_321_14 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_321_15 <= 1'h0;
    end else begin
      if (_T_382) begin
        if (4'hf == io_in_0_d_bits_source) begin
          _T_321_15 <= 1'h0;
        end else begin
          if (_T_375) begin
            if (4'hf == io_in_0_a_bits_source) begin
              _T_321_15 <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_375) begin
          if (4'hf == io_in_0_a_bits_source) begin
            _T_321_15 <= 1'h1;
          end
        end
      end
    end
    if (_T_400) begin
      _T_405 <= _T_182;
    end
    if (_T_431) begin
      _T_436 <= _T_182;
    end
  end
endmodule
module TLXbar_1(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_4_a_ready,
  output        io_out_4_a_valid,
  output [2:0]  io_out_4_a_bits_opcode,
  output [2:0]  io_out_4_a_bits_param,
  output [2:0]  io_out_4_a_bits_size,
  output [4:0]  io_out_4_a_bits_source,
  output [31:0] io_out_4_a_bits_address,
  output [3:0]  io_out_4_a_bits_mask,
  output [31:0] io_out_4_a_bits_data,
  output        io_out_4_d_ready,
  input         io_out_4_d_valid,
  input  [2:0]  io_out_4_d_bits_opcode,
  input  [1:0]  io_out_4_d_bits_param,
  input  [2:0]  io_out_4_d_bits_size,
  input  [4:0]  io_out_4_d_bits_source,
  input         io_out_4_d_bits_sink,
  input  [31:0] io_out_4_d_bits_data,
  input         io_out_4_d_bits_error,
  input         io_out_3_a_ready,
  output        io_out_3_a_valid,
  output [2:0]  io_out_3_a_bits_opcode,
  output [2:0]  io_out_3_a_bits_size,
  output [4:0]  io_out_3_a_bits_source,
  output [16:0] io_out_3_a_bits_address,
  output [3:0]  io_out_3_a_bits_mask,
  output        io_out_3_d_ready,
  input         io_out_3_d_valid,
  input  [2:0]  io_out_3_d_bits_opcode,
  input  [1:0]  io_out_3_d_bits_param,
  input  [2:0]  io_out_3_d_bits_size,
  input  [4:0]  io_out_3_d_bits_source,
  input         io_out_3_d_bits_sink,
  input  [31:0] io_out_3_d_bits_data,
  input         io_out_3_d_bits_error,
  input         io_out_2_a_ready,
  output        io_out_2_a_valid,
  output [2:0]  io_out_2_a_bits_opcode,
  output [2:0]  io_out_2_a_bits_size,
  output [4:0]  io_out_2_a_bits_source,
  output [11:0] io_out_2_a_bits_address,
  output [3:0]  io_out_2_a_bits_mask,
  output [31:0] io_out_2_a_bits_data,
  output        io_out_2_d_ready,
  input         io_out_2_d_valid,
  input  [2:0]  io_out_2_d_bits_opcode,
  input  [1:0]  io_out_2_d_bits_param,
  input  [2:0]  io_out_2_d_bits_size,
  input  [4:0]  io_out_2_d_bits_source,
  input         io_out_2_d_bits_sink,
  input  [31:0] io_out_2_d_bits_data,
  input         io_out_2_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [2:0]  io_out_1_a_bits_size,
  output [4:0]  io_out_1_a_bits_source,
  output [25:0] io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [2:0]  io_out_1_d_bits_size,
  input  [4:0]  io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [31:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [27:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire [31:0] _T_1000;
  wire [32:0] _T_1001;
  wire [32:0] _T_1003;
  wire [32:0] _T_1004;
  wire  _T_1006;
  wire [31:0] _T_1008;
  wire [32:0] _T_1009;
  wire [32:0] _T_1011;
  wire [32:0] _T_1012;
  wire  _T_1014;
  wire [32:0] _T_1017;
  wire [32:0] _T_1019;
  wire [32:0] _T_1020;
  wire  _T_1022;
  wire [31:0] _T_1024;
  wire [32:0] _T_1025;
  wire [32:0] _T_1027;
  wire [32:0] _T_1028;
  wire  _T_1030;
  wire [31:0] _T_1032;
  wire [32:0] _T_1033;
  wire [32:0] _T_1035;
  wire [32:0] _T_1036;
  wire  _T_1038;
  wire [12:0] _T_1903;
  wire [5:0] _T_1904;
  wire [5:0] _T_1905;
  wire [3:0] _T_1906;
  wire  _T_1907;
  wire [3:0] _T_1909;
  wire [12:0] _T_1912;
  wire [5:0] _T_1913;
  wire [5:0] _T_1914;
  wire [3:0] _T_1915;
  wire  _T_1916;
  wire [3:0] _T_1918;
  wire [12:0] _T_1921;
  wire [5:0] _T_1922;
  wire [5:0] _T_1923;
  wire [3:0] _T_1924;
  wire  _T_1925;
  wire [3:0] _T_1927;
  wire [12:0] _T_1930;
  wire [5:0] _T_1931;
  wire [5:0] _T_1932;
  wire [3:0] _T_1933;
  wire [12:0] _T_1940;
  wire [5:0] _T_1941;
  wire [5:0] _T_1942;
  wire [3:0] _T_1943;
  wire  _T_1944;
  wire [3:0] _T_1946;
  wire  _T_2026;
  wire  _T_2027;
  wire  _T_2028;
  wire  _T_2029;
  wire  _T_2030;
  wire  _T_2033;
  wire  _T_2035;
  wire  _T_2037;
  wire  _T_2039;
  wire  _T_2041;
  wire  _T_2042;
  wire  _T_2043;
  wire  _T_2044;
  wire  _T_2045;
  wire  _T_2496;
  wire  _T_2503;
  wire  _T_2504;
  wire  _T_2506;
  wire  _T_2570;
  wire  _T_2577;
  wire  _T_2578;
  wire  _T_2580;
  wire  _T_2644;
  wire  _T_2651;
  wire  _T_2652;
  wire  _T_2654;
  wire  _T_2718;
  wire  _T_2725;
  wire  _T_2726;
  wire  _T_2728;
  wire  _T_2792;
  wire  _T_2799;
  wire  _T_2800;
  wire  _T_2802;
  reg [3:0] _T_2843;
  reg [31:0] _RAND_0;
  wire  _T_2845;
  wire  _T_2846;
  wire [1:0] _T_2847;
  wire [1:0] _T_2848;
  wire [2:0] _T_2849;
  wire [4:0] _T_2850;
  wire  _T_2852;
  wire  _T_2853;
  wire  _T_2855;
  reg [4:0] _T_2859;
  reg [31:0] _RAND_1;
  wire [4:0] _T_2860;
  wire [4:0] _T_2861;
  wire [9:0] _T_2862;
  wire [8:0] _T_2863;
  wire [9:0] _GEN_6;
  wire [9:0] _T_2864;
  wire [7:0] _T_2865;
  wire [9:0] _GEN_7;
  wire [9:0] _T_2866;
  wire [5:0] _T_2867;
  wire [9:0] _GEN_8;
  wire [9:0] _T_2868;
  wire [8:0] _T_2870;
  wire [9:0] _GEN_9;
  wire [9:0] _T_2871;
  wire [9:0] _GEN_10;
  wire [9:0] _T_2872;
  wire [4:0] _T_2873;
  wire [4:0] _T_2874;
  wire [4:0] _T_2875;
  wire [4:0] _T_2876;
  wire  _T_2878;
  wire  _T_2879;
  wire [4:0] _T_2880;
  wire [5:0] _GEN_11;
  wire [5:0] _T_2881;
  wire [4:0] _T_2882;
  wire [4:0] _T_2883;
  wire [6:0] _GEN_12;
  wire [6:0] _T_2884;
  wire [4:0] _T_2885;
  wire [4:0] _T_2886;
  wire [8:0] _GEN_13;
  wire [8:0] _T_2887;
  wire [4:0] _T_2888;
  wire [4:0] _T_2889;
  wire [4:0] _GEN_0;
  wire  _T_2892;
  wire  _T_2893;
  wire  _T_2894;
  wire  _T_2895;
  wire  _T_2896;
  wire  _T_2907;
  wire  _T_2908;
  wire  _T_2909;
  wire  _T_2910;
  wire  _T_2911;
  wire  _T_2924;
  wire  _T_2925;
  wire  _T_2926;
  wire  _T_2927;
  wire  _T_2931;
  wire  _T_2936;
  wire  _T_2937;
  wire  _T_2939;
  wire  _T_2941;
  wire  _T_2942;
  wire  _T_2944;
  wire  _T_2946;
  wire  _T_2947;
  wire  _T_2949;
  wire  _T_2951;
  wire  _T_2952;
  wire  _T_2954;
  wire  _T_2955;
  wire  _T_2956;
  wire  _T_2957;
  wire  _T_2959;
  wire  _T_2960;
  wire  _T_2961;
  wire  _T_2962;
  wire  _T_2963;
  wire  _T_2965;
  wire  _T_2970;
  wire  _T_2971;
  wire  _T_2973;
  wire [3:0] _T_2975;
  wire [3:0] _T_2977;
  wire [3:0] _T_2979;
  wire [3:0] _T_2981;
  wire [3:0] _T_2983;
  wire [3:0] _T_2984;
  wire [3:0] _T_2985;
  wire [3:0] _T_2986;
  wire [3:0] _T_2987;
  wire  _T_2988;
  wire [3:0] _GEN_14;
  wire [4:0] _T_2989;
  wire [4:0] _T_2990;
  wire [3:0] _T_2991;
  wire [3:0] _T_2992;
  reg  _T_3022_0;
  reg [31:0] _RAND_2;
  reg  _T_3022_1;
  reg [31:0] _RAND_3;
  reg  _T_3022_2;
  reg [31:0] _RAND_4;
  reg  _T_3022_3;
  reg [31:0] _RAND_5;
  reg  _T_3022_4;
  reg [31:0] _RAND_6;
  wire  _T_3042_0;
  wire  _T_3042_1;
  wire  _T_3042_2;
  wire  _T_3042_3;
  wire  _T_3042_4;
  wire  _T_3056_0;
  wire  _T_3056_1;
  wire  _T_3056_2;
  wire  _T_3056_3;
  wire  _T_3056_4;
  wire  _T_3070;
  wire  _T_3071;
  wire  _T_3072;
  wire  _T_3073;
  wire  _T_3074;
  wire  _T_3081;
  wire  _T_3083;
  wire  _T_3085;
  wire  _T_3087;
  wire  _T_3089;
  wire  _T_3090;
  wire  _T_3091;
  wire  _T_3092;
  wire  _T_3093;
  wire  _T_3096;
  wire [32:0] _T_3098;
  wire [33:0] _T_3099;
  wire [7:0] _T_3100;
  wire [4:0] _T_3101;
  wire [12:0] _T_3102;
  wire [46:0] _T_3103;
  wire [46:0] _T_3105;
  wire [32:0] _T_3106;
  wire [33:0] _T_3107;
  wire [7:0] _T_3108;
  wire [4:0] _T_3109;
  wire [12:0] _T_3110;
  wire [46:0] _T_3111;
  wire [46:0] _T_3113;
  wire [32:0] _T_3114;
  wire [33:0] _T_3115;
  wire [7:0] _T_3116;
  wire [4:0] _T_3117;
  wire [12:0] _T_3118;
  wire [46:0] _T_3119;
  wire [46:0] _T_3121;
  wire [32:0] _T_3122;
  wire [33:0] _T_3123;
  wire [7:0] _T_3124;
  wire [4:0] _T_3125;
  wire [12:0] _T_3126;
  wire [46:0] _T_3127;
  wire [46:0] _T_3129;
  wire [32:0] _T_3130;
  wire [33:0] _T_3131;
  wire [7:0] _T_3132;
  wire [4:0] _T_3133;
  wire [12:0] _T_3134;
  wire [46:0] _T_3135;
  wire [46:0] _T_3137;
  wire [46:0] _T_3138;
  wire [46:0] _T_3139;
  wire [46:0] _T_3140;
  wire [46:0] _T_3141;
  wire  _T_3146;
  wire [31:0] _T_3147;
  wire  _T_3148;
  wire [4:0] _T_3149;
  wire [2:0] _T_3150;
  wire [1:0] _T_3151;
  wire [2:0] _T_3152;
  assign io_in_0_a_ready = _T_2045;
  assign io_in_0_d_valid = _T_3096;
  assign io_in_0_d_bits_opcode = _T_3152;
  assign io_in_0_d_bits_param = _T_3151;
  assign io_in_0_d_bits_size = _T_3150;
  assign io_in_0_d_bits_source = _T_3149;
  assign io_in_0_d_bits_sink = _T_3148;
  assign io_in_0_d_bits_data = _T_3147;
  assign io_in_0_d_bits_error = _T_3146;
  assign io_out_4_a_valid = _T_2030;
  assign io_out_4_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_4_a_bits_param = io_in_0_a_bits_param;
  assign io_out_4_a_bits_size = io_in_0_a_bits_size;
  assign io_out_4_a_bits_source = io_in_0_a_bits_source;
  assign io_out_4_a_bits_address = io_in_0_a_bits_address;
  assign io_out_4_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_4_a_bits_data = io_in_0_a_bits_data;
  assign io_out_4_d_ready = _T_3074;
  assign io_out_3_a_valid = _T_2029;
  assign io_out_3_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_3_a_bits_size = io_in_0_a_bits_size;
  assign io_out_3_a_bits_source = io_in_0_a_bits_source;
  assign io_out_3_a_bits_address = io_in_0_a_bits_address[16:0];
  assign io_out_3_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_3_d_ready = _T_3073;
  assign io_out_2_a_valid = _T_2028;
  assign io_out_2_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_2_a_bits_size = io_in_0_a_bits_size;
  assign io_out_2_a_bits_source = io_in_0_a_bits_source;
  assign io_out_2_a_bits_address = io_in_0_a_bits_address[11:0];
  assign io_out_2_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_2_a_bits_data = io_in_0_a_bits_data;
  assign io_out_2_d_ready = _T_3072;
  assign io_out_1_a_valid = _T_2027;
  assign io_out_1_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_1_a_bits_size = io_in_0_a_bits_size;
  assign io_out_1_a_bits_source = io_in_0_a_bits_source;
  assign io_out_1_a_bits_address = io_in_0_a_bits_address[25:0];
  assign io_out_1_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_1_a_bits_data = io_in_0_a_bits_data;
  assign io_out_1_d_ready = _T_3071;
  assign io_out_0_a_valid = _T_2026;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address[27:0];
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = _T_3070;
  assign _T_1000 = io_in_0_a_bits_address ^ 32'h4000000;
  assign _T_1001 = {1'b0,$signed(_T_1000)};
  assign _T_1003 = $signed(_T_1001) & $signed(33'sh84000000);
  assign _T_1004 = $signed(_T_1003);
  assign _T_1006 = $signed(_T_1004) == $signed(33'sh0);
  assign _T_1008 = io_in_0_a_bits_address ^ 32'h2000000;
  assign _T_1009 = {1'b0,$signed(_T_1008)};
  assign _T_1011 = $signed(_T_1009) & $signed(33'sh86010000);
  assign _T_1012 = $signed(_T_1011);
  assign _T_1014 = $signed(_T_1012) == $signed(33'sh0);
  assign _T_1017 = {1'b0,$signed(io_in_0_a_bits_address)};
  assign _T_1019 = $signed(_T_1017) & $signed(33'sh86010000);
  assign _T_1020 = $signed(_T_1019);
  assign _T_1022 = $signed(_T_1020) == $signed(33'sh0);
  assign _T_1024 = io_in_0_a_bits_address ^ 32'h10000;
  assign _T_1025 = {1'b0,$signed(_T_1024)};
  assign _T_1027 = $signed(_T_1025) & $signed(33'sh86010000);
  assign _T_1028 = $signed(_T_1027);
  assign _T_1030 = $signed(_T_1028) == $signed(33'sh0);
  assign _T_1032 = io_in_0_a_bits_address ^ 32'h80000000;
  assign _T_1033 = {1'b0,$signed(_T_1032)};
  assign _T_1035 = $signed(_T_1033) & $signed(33'sh86010000);
  assign _T_1036 = $signed(_T_1035);
  assign _T_1038 = $signed(_T_1036) == $signed(33'sh0);
  assign _T_1903 = 13'h3f << io_out_0_d_bits_size;
  assign _T_1904 = _T_1903[5:0];
  assign _T_1905 = ~ _T_1904;
  assign _T_1906 = _T_1905[5:2];
  assign _T_1907 = io_out_0_d_bits_opcode[0];
  assign _T_1909 = _T_1907 ? _T_1906 : 4'h0;
  assign _T_1912 = 13'h3f << io_out_1_d_bits_size;
  assign _T_1913 = _T_1912[5:0];
  assign _T_1914 = ~ _T_1913;
  assign _T_1915 = _T_1914[5:2];
  assign _T_1916 = io_out_1_d_bits_opcode[0];
  assign _T_1918 = _T_1916 ? _T_1915 : 4'h0;
  assign _T_1921 = 13'h3f << io_out_2_d_bits_size;
  assign _T_1922 = _T_1921[5:0];
  assign _T_1923 = ~ _T_1922;
  assign _T_1924 = _T_1923[5:2];
  assign _T_1925 = io_out_2_d_bits_opcode[0];
  assign _T_1927 = _T_1925 ? _T_1924 : 4'h0;
  assign _T_1930 = 13'h3f << io_out_3_d_bits_size;
  assign _T_1931 = _T_1930[5:0];
  assign _T_1932 = ~ _T_1931;
  assign _T_1933 = _T_1932[5:2];
  assign _T_1940 = 13'h3f << io_out_4_d_bits_size;
  assign _T_1941 = _T_1940[5:0];
  assign _T_1942 = ~ _T_1941;
  assign _T_1943 = _T_1942[5:2];
  assign _T_1944 = io_out_4_d_bits_opcode[0];
  assign _T_1946 = _T_1944 ? _T_1943 : 4'h0;
  assign _T_2026 = io_in_0_a_valid & _T_1006;
  assign _T_2027 = io_in_0_a_valid & _T_1014;
  assign _T_2028 = io_in_0_a_valid & _T_1022;
  assign _T_2029 = io_in_0_a_valid & _T_1030;
  assign _T_2030 = io_in_0_a_valid & _T_1038;
  assign _T_2033 = _T_1006 ? io_out_0_a_ready : 1'h0;
  assign _T_2035 = _T_1014 ? io_out_1_a_ready : 1'h0;
  assign _T_2037 = _T_1022 ? io_out_2_a_ready : 1'h0;
  assign _T_2039 = _T_1030 ? io_out_3_a_ready : 1'h0;
  assign _T_2041 = _T_1038 ? io_out_4_a_ready : 1'h0;
  assign _T_2042 = _T_2033 | _T_2035;
  assign _T_2043 = _T_2042 | _T_2037;
  assign _T_2044 = _T_2043 | _T_2039;
  assign _T_2045 = _T_2044 | _T_2041;
  assign _T_2496 = _T_2026 == 1'h0;
  assign _T_2503 = _T_2496 | _T_2026;
  assign _T_2504 = _T_2503 | reset;
  assign _T_2506 = _T_2504 == 1'h0;
  assign _T_2570 = _T_2027 == 1'h0;
  assign _T_2577 = _T_2570 | _T_2027;
  assign _T_2578 = _T_2577 | reset;
  assign _T_2580 = _T_2578 == 1'h0;
  assign _T_2644 = _T_2028 == 1'h0;
  assign _T_2651 = _T_2644 | _T_2028;
  assign _T_2652 = _T_2651 | reset;
  assign _T_2654 = _T_2652 == 1'h0;
  assign _T_2718 = _T_2029 == 1'h0;
  assign _T_2725 = _T_2718 | _T_2029;
  assign _T_2726 = _T_2725 | reset;
  assign _T_2728 = _T_2726 == 1'h0;
  assign _T_2792 = _T_2030 == 1'h0;
  assign _T_2799 = _T_2792 | _T_2030;
  assign _T_2800 = _T_2799 | reset;
  assign _T_2802 = _T_2800 == 1'h0;
  assign _T_2845 = _T_2843 == 4'h0;
  assign _T_2846 = _T_2845 & io_in_0_d_ready;
  assign _T_2847 = {io_out_1_d_valid,io_out_0_d_valid};
  assign _T_2848 = {io_out_4_d_valid,io_out_3_d_valid};
  assign _T_2849 = {_T_2848,io_out_2_d_valid};
  assign _T_2850 = {_T_2849,_T_2847};
  assign _T_2852 = _T_2850 == _T_2850;
  assign _T_2853 = _T_2852 | reset;
  assign _T_2855 = _T_2853 == 1'h0;
  assign _T_2860 = ~ _T_2859;
  assign _T_2861 = _T_2850 & _T_2860;
  assign _T_2862 = {_T_2861,_T_2850};
  assign _T_2863 = _T_2862[9:1];
  assign _GEN_6 = {{1'd0}, _T_2863};
  assign _T_2864 = _T_2862 | _GEN_6;
  assign _T_2865 = _T_2864[9:2];
  assign _GEN_7 = {{2'd0}, _T_2865};
  assign _T_2866 = _T_2864 | _GEN_7;
  assign _T_2867 = _T_2866[9:4];
  assign _GEN_8 = {{4'd0}, _T_2867};
  assign _T_2868 = _T_2866 | _GEN_8;
  assign _T_2870 = _T_2868[9:1];
  assign _GEN_9 = {{5'd0}, _T_2859};
  assign _T_2871 = _GEN_9 << 5;
  assign _GEN_10 = {{1'd0}, _T_2870};
  assign _T_2872 = _GEN_10 | _T_2871;
  assign _T_2873 = _T_2872[9:5];
  assign _T_2874 = _T_2872[4:0];
  assign _T_2875 = _T_2873 & _T_2874;
  assign _T_2876 = ~ _T_2875;
  assign _T_2878 = _T_2850 != 5'h0;
  assign _T_2879 = _T_2846 & _T_2878;
  assign _T_2880 = _T_2876 & _T_2850;
  assign _GEN_11 = {{1'd0}, _T_2880};
  assign _T_2881 = _GEN_11 << 1;
  assign _T_2882 = _T_2881[4:0];
  assign _T_2883 = _T_2880 | _T_2882;
  assign _GEN_12 = {{2'd0}, _T_2883};
  assign _T_2884 = _GEN_12 << 2;
  assign _T_2885 = _T_2884[4:0];
  assign _T_2886 = _T_2883 | _T_2885;
  assign _GEN_13 = {{4'd0}, _T_2886};
  assign _T_2887 = _GEN_13 << 4;
  assign _T_2888 = _T_2887[4:0];
  assign _T_2889 = _T_2886 | _T_2888;
  assign _GEN_0 = _T_2879 ? _T_2889 : _T_2859;
  assign _T_2892 = _T_2876[0];
  assign _T_2893 = _T_2876[1];
  assign _T_2894 = _T_2876[2];
  assign _T_2895 = _T_2876[3];
  assign _T_2896 = _T_2876[4];
  assign _T_2907 = _T_2892 & io_out_0_d_valid;
  assign _T_2908 = _T_2893 & io_out_1_d_valid;
  assign _T_2909 = _T_2894 & io_out_2_d_valid;
  assign _T_2910 = _T_2895 & io_out_3_d_valid;
  assign _T_2911 = _T_2896 & io_out_4_d_valid;
  assign _T_2924 = _T_2907 | _T_2908;
  assign _T_2925 = _T_2924 | _T_2909;
  assign _T_2926 = _T_2925 | _T_2910;
  assign _T_2927 = _T_2926 | _T_2911;
  assign _T_2931 = _T_2907 == 1'h0;
  assign _T_2936 = _T_2908 == 1'h0;
  assign _T_2937 = _T_2931 | _T_2936;
  assign _T_2939 = _T_2924 == 1'h0;
  assign _T_2941 = _T_2909 == 1'h0;
  assign _T_2942 = _T_2939 | _T_2941;
  assign _T_2944 = _T_2925 == 1'h0;
  assign _T_2946 = _T_2910 == 1'h0;
  assign _T_2947 = _T_2944 | _T_2946;
  assign _T_2949 = _T_2926 == 1'h0;
  assign _T_2951 = _T_2911 == 1'h0;
  assign _T_2952 = _T_2949 | _T_2951;
  assign _T_2954 = _T_2937 & _T_2942;
  assign _T_2955 = _T_2954 & _T_2947;
  assign _T_2956 = _T_2955 & _T_2952;
  assign _T_2957 = _T_2956 | reset;
  assign _T_2959 = _T_2957 == 1'h0;
  assign _T_2960 = io_out_0_d_valid | io_out_1_d_valid;
  assign _T_2961 = _T_2960 | io_out_2_d_valid;
  assign _T_2962 = _T_2961 | io_out_3_d_valid;
  assign _T_2963 = _T_2962 | io_out_4_d_valid;
  assign _T_2965 = _T_2963 == 1'h0;
  assign _T_2970 = _T_2965 | _T_2927;
  assign _T_2971 = _T_2970 | reset;
  assign _T_2973 = _T_2971 == 1'h0;
  assign _T_2975 = _T_2907 ? _T_1909 : 4'h0;
  assign _T_2977 = _T_2908 ? _T_1918 : 4'h0;
  assign _T_2979 = _T_2909 ? _T_1927 : 4'h0;
  assign _T_2981 = _T_2910 ? _T_1933 : 4'h0;
  assign _T_2983 = _T_2911 ? _T_1946 : 4'h0;
  assign _T_2984 = _T_2975 | _T_2977;
  assign _T_2985 = _T_2984 | _T_2979;
  assign _T_2986 = _T_2985 | _T_2981;
  assign _T_2987 = _T_2986 | _T_2983;
  assign _T_2988 = io_in_0_d_ready & _T_3096;
  assign _GEN_14 = {{3'd0}, _T_2988};
  assign _T_2989 = _T_2843 - _GEN_14;
  assign _T_2990 = $unsigned(_T_2989);
  assign _T_2991 = _T_2990[3:0];
  assign _T_2992 = _T_2846 ? _T_2987 : _T_2991;
  assign _T_3042_0 = _T_2845 ? _T_2907 : _T_3022_0;
  assign _T_3042_1 = _T_2845 ? _T_2908 : _T_3022_1;
  assign _T_3042_2 = _T_2845 ? _T_2909 : _T_3022_2;
  assign _T_3042_3 = _T_2845 ? _T_2910 : _T_3022_3;
  assign _T_3042_4 = _T_2845 ? _T_2911 : _T_3022_4;
  assign _T_3056_0 = _T_2845 ? _T_2892 : _T_3022_0;
  assign _T_3056_1 = _T_2845 ? _T_2893 : _T_3022_1;
  assign _T_3056_2 = _T_2845 ? _T_2894 : _T_3022_2;
  assign _T_3056_3 = _T_2845 ? _T_2895 : _T_3022_3;
  assign _T_3056_4 = _T_2845 ? _T_2896 : _T_3022_4;
  assign _T_3070 = io_in_0_d_ready & _T_3056_0;
  assign _T_3071 = io_in_0_d_ready & _T_3056_1;
  assign _T_3072 = io_in_0_d_ready & _T_3056_2;
  assign _T_3073 = io_in_0_d_ready & _T_3056_3;
  assign _T_3074 = io_in_0_d_ready & _T_3056_4;
  assign _T_3081 = _T_3022_0 ? io_out_0_d_valid : 1'h0;
  assign _T_3083 = _T_3022_1 ? io_out_1_d_valid : 1'h0;
  assign _T_3085 = _T_3022_2 ? io_out_2_d_valid : 1'h0;
  assign _T_3087 = _T_3022_3 ? io_out_3_d_valid : 1'h0;
  assign _T_3089 = _T_3022_4 ? io_out_4_d_valid : 1'h0;
  assign _T_3090 = _T_3081 | _T_3083;
  assign _T_3091 = _T_3090 | _T_3085;
  assign _T_3092 = _T_3091 | _T_3087;
  assign _T_3093 = _T_3092 | _T_3089;
  assign _T_3096 = _T_2845 ? _T_2963 : _T_3093;
  assign _T_3098 = {io_out_0_d_bits_sink,io_out_0_d_bits_data};
  assign _T_3099 = {_T_3098,io_out_0_d_bits_error};
  assign _T_3100 = {io_out_0_d_bits_size,io_out_0_d_bits_source};
  assign _T_3101 = {io_out_0_d_bits_opcode,io_out_0_d_bits_param};
  assign _T_3102 = {_T_3101,_T_3100};
  assign _T_3103 = {_T_3102,_T_3099};
  assign _T_3105 = _T_3042_0 ? _T_3103 : 47'h0;
  assign _T_3106 = {io_out_1_d_bits_sink,io_out_1_d_bits_data};
  assign _T_3107 = {_T_3106,io_out_1_d_bits_error};
  assign _T_3108 = {io_out_1_d_bits_size,io_out_1_d_bits_source};
  assign _T_3109 = {io_out_1_d_bits_opcode,io_out_1_d_bits_param};
  assign _T_3110 = {_T_3109,_T_3108};
  assign _T_3111 = {_T_3110,_T_3107};
  assign _T_3113 = _T_3042_1 ? _T_3111 : 47'h0;
  assign _T_3114 = {io_out_2_d_bits_sink,io_out_2_d_bits_data};
  assign _T_3115 = {_T_3114,io_out_2_d_bits_error};
  assign _T_3116 = {io_out_2_d_bits_size,io_out_2_d_bits_source};
  assign _T_3117 = {io_out_2_d_bits_opcode,io_out_2_d_bits_param};
  assign _T_3118 = {_T_3117,_T_3116};
  assign _T_3119 = {_T_3118,_T_3115};
  assign _T_3121 = _T_3042_2 ? _T_3119 : 47'h0;
  assign _T_3122 = {io_out_3_d_bits_sink,io_out_3_d_bits_data};
  assign _T_3123 = {_T_3122,io_out_3_d_bits_error};
  assign _T_3124 = {io_out_3_d_bits_size,io_out_3_d_bits_source};
  assign _T_3125 = {io_out_3_d_bits_opcode,io_out_3_d_bits_param};
  assign _T_3126 = {_T_3125,_T_3124};
  assign _T_3127 = {_T_3126,_T_3123};
  assign _T_3129 = _T_3042_3 ? _T_3127 : 47'h0;
  assign _T_3130 = {io_out_4_d_bits_sink,io_out_4_d_bits_data};
  assign _T_3131 = {_T_3130,io_out_4_d_bits_error};
  assign _T_3132 = {io_out_4_d_bits_size,io_out_4_d_bits_source};
  assign _T_3133 = {io_out_4_d_bits_opcode,io_out_4_d_bits_param};
  assign _T_3134 = {_T_3133,_T_3132};
  assign _T_3135 = {_T_3134,_T_3131};
  assign _T_3137 = _T_3042_4 ? _T_3135 : 47'h0;
  assign _T_3138 = _T_3105 | _T_3113;
  assign _T_3139 = _T_3138 | _T_3121;
  assign _T_3140 = _T_3139 | _T_3129;
  assign _T_3141 = _T_3140 | _T_3137;
  assign _T_3146 = _T_3141[0];
  assign _T_3147 = _T_3141[32:1];
  assign _T_3148 = _T_3141[33];
  assign _T_3149 = _T_3141[38:34];
  assign _T_3150 = _T_3141[41:39];
  assign _T_3151 = _T_3141[43:42];
  assign _T_3152 = _T_3141[46:44];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_2843 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_2859 = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_3022_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_3022_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_3022_2 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_3022_3 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_3022_4 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_2843 <= 4'h0;
    end else begin
      if (_T_2846) begin
        _T_2843 <= _T_2987;
      end else begin
        _T_2843 <= _T_2991;
      end
    end
    if (reset) begin
      _T_2859 <= 5'h1f;
    end else begin
      if (_T_2879) begin
        _T_2859 <= _T_2889;
      end
    end
    if (reset) begin
      _T_3022_0 <= 1'h0;
    end else begin
      if (_T_2845) begin
        _T_3022_0 <= _T_2907;
      end
    end
    if (reset) begin
      _T_3022_1 <= 1'h0;
    end else begin
      if (_T_2845) begin
        _T_3022_1 <= _T_2908;
      end
    end
    if (reset) begin
      _T_3022_2 <= 1'h0;
    end else begin
      if (_T_2845) begin
        _T_3022_2 <= _T_2909;
      end
    end
    if (reset) begin
      _T_3022_3 <= 1'h0;
    end else begin
      if (_T_2845) begin
        _T_3022_3 <= _T_2910;
      end
    end
    if (reset) begin
      _T_3022_4 <= 1'h0;
    end else begin
      if (_T_2845) begin
        _T_3022_4 <= _T_2911;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2506) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2506) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2580) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2654) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2654) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2728) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2728) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2802) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2802) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2855) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2855) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2959) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2959) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2973) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2973) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_6(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_43_data;
  wire  ram_opcode__T_43_addr;
  wire [2:0] ram_opcode__T_29_data;
  wire  ram_opcode__T_29_addr;
  wire  ram_opcode__T_29_mask;
  wire  ram_opcode__T_29_en;
  reg [2:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_43_data;
  wire  ram_param__T_43_addr;
  wire [2:0] ram_param__T_29_data;
  wire  ram_param__T_29_addr;
  wire  ram_param__T_29_mask;
  wire  ram_param__T_29_en;
  reg [2:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [2:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [2:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg [4:0] ram_source [0:1];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_43_data;
  wire  ram_source__T_43_addr;
  wire [4:0] ram_source__T_29_data;
  wire  ram_source__T_29_addr;
  wire  ram_source__T_29_mask;
  wire  ram_source__T_29_en;
  reg [31:0] ram_address [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_43_data;
  wire  ram_address__T_43_addr;
  wire [31:0] ram_address__T_29_data;
  wire  ram_address__T_29_addr;
  wire  ram_address__T_29_mask;
  wire  ram_address__T_29_en;
  reg [3:0] ram_mask [0:1];
  reg [31:0] _RAND_5;
  wire [3:0] ram_mask__T_43_data;
  wire  ram_mask__T_43_addr;
  wire [3:0] ram_mask__T_29_data;
  wire  ram_mask__T_29_addr;
  wire  ram_mask__T_29_mask;
  wire  ram_mask__T_29_en;
  reg [31:0] ram_data [0:1];
  reg [31:0] _RAND_6;
  wire [31:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [31:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg  value;
  reg [31:0] _RAND_7;
  reg  value_1;
  reg [31:0] _RAND_8;
  reg  maybe_full;
  reg [31:0] _RAND_9;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_10;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_11;
  wire  _T_38;
  wire  _GEN_12;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_opcode = ram_opcode__T_43_data;
  assign io_deq_bits_param = ram_param__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_source = ram_source__T_43_data;
  assign io_deq_bits_address = ram_address__T_43_data;
  assign io_deq_bits_mask = ram_mask__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign ram_opcode__T_43_addr = value_1;
  assign ram_opcode__T_43_data = ram_opcode[ram_opcode__T_43_addr];
  assign ram_opcode__T_29_data = io_enq_bits_opcode;
  assign ram_opcode__T_29_addr = value;
  assign ram_opcode__T_29_mask = _T_25;
  assign ram_opcode__T_29_en = _T_25;
  assign ram_param__T_43_addr = value_1;
  assign ram_param__T_43_data = ram_param[ram_param__T_43_addr];
  assign ram_param__T_29_data = io_enq_bits_param;
  assign ram_param__T_29_addr = value;
  assign ram_param__T_29_mask = _T_25;
  assign ram_param__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_source__T_43_addr = value_1;
  assign ram_source__T_43_data = ram_source[ram_source__T_43_addr];
  assign ram_source__T_29_data = io_enq_bits_source;
  assign ram_source__T_29_addr = value;
  assign ram_source__T_29_mask = _T_25;
  assign ram_source__T_29_en = _T_25;
  assign ram_address__T_43_addr = value_1;
  assign ram_address__T_43_data = ram_address[ram_address__T_43_addr];
  assign ram_address__T_29_data = io_enq_bits_address;
  assign ram_address__T_29_addr = value;
  assign ram_address__T_29_mask = _T_25;
  assign ram_address__T_29_en = _T_25;
  assign ram_mask__T_43_addr = value_1;
  assign ram_mask__T_43_data = ram_mask[ram_mask__T_43_addr];
  assign ram_mask__T_29_data = io_enq_bits_mask;
  assign ram_mask__T_29_addr = value;
  assign ram_mask__T_29_mask = _T_25;
  assign ram_mask__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_10 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_11 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_12 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_29_en & ram_opcode__T_29_mask) begin
      ram_opcode[ram_opcode__T_29_addr] <= ram_opcode__T_29_data;
    end
    if(ram_param__T_29_en & ram_param__T_29_mask) begin
      ram_param[ram_param__T_29_addr] <= ram_param__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_source__T_29_en & ram_source__T_29_mask) begin
      ram_source[ram_source__T_29_addr] <= ram_source__T_29_data;
    end
    if(ram_address__T_29_en & ram_address__T_29_mask) begin
      ram_address[ram_address__T_29_addr] <= ram_address__T_29_data;
    end
    if(ram_mask__T_29_en & ram_mask__T_29_mask) begin
      ram_mask[ram_mask__T_29_addr] <= ram_mask__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_7(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input         io_enq_bits_sink,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output        io_deq_bits_sink,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_43_data;
  wire  ram_opcode__T_43_addr;
  wire [2:0] ram_opcode__T_29_data;
  wire  ram_opcode__T_29_addr;
  wire  ram_opcode__T_29_mask;
  wire  ram_opcode__T_29_en;
  reg [1:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_43_data;
  wire  ram_param__T_43_addr;
  wire [1:0] ram_param__T_29_data;
  wire  ram_param__T_29_addr;
  wire  ram_param__T_29_mask;
  wire  ram_param__T_29_en;
  reg [2:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [2:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [2:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg [4:0] ram_source [0:1];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_43_data;
  wire  ram_source__T_43_addr;
  wire [4:0] ram_source__T_29_data;
  wire  ram_source__T_29_addr;
  wire  ram_source__T_29_mask;
  wire  ram_source__T_29_en;
  reg  ram_sink [0:1];
  reg [31:0] _RAND_4;
  wire  ram_sink__T_43_data;
  wire  ram_sink__T_43_addr;
  wire  ram_sink__T_29_data;
  wire  ram_sink__T_29_addr;
  wire  ram_sink__T_29_mask;
  wire  ram_sink__T_29_en;
  reg [31:0] ram_data [0:1];
  reg [31:0] _RAND_5;
  wire [31:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [31:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg  ram_error [0:1];
  reg [31:0] _RAND_6;
  wire  ram_error__T_43_data;
  wire  ram_error__T_43_addr;
  wire  ram_error__T_29_data;
  wire  ram_error__T_29_addr;
  wire  ram_error__T_29_mask;
  wire  ram_error__T_29_en;
  reg  value;
  reg [31:0] _RAND_7;
  reg  value_1;
  reg [31:0] _RAND_8;
  reg  maybe_full;
  reg [31:0] _RAND_9;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_10;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_11;
  wire  _T_38;
  wire  _GEN_12;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_opcode = ram_opcode__T_43_data;
  assign io_deq_bits_param = ram_param__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_source = ram_source__T_43_data;
  assign io_deq_bits_sink = ram_sink__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign io_deq_bits_error = ram_error__T_43_data;
  assign ram_opcode__T_43_addr = value_1;
  assign ram_opcode__T_43_data = ram_opcode[ram_opcode__T_43_addr];
  assign ram_opcode__T_29_data = io_enq_bits_opcode;
  assign ram_opcode__T_29_addr = value;
  assign ram_opcode__T_29_mask = _T_25;
  assign ram_opcode__T_29_en = _T_25;
  assign ram_param__T_43_addr = value_1;
  assign ram_param__T_43_data = ram_param[ram_param__T_43_addr];
  assign ram_param__T_29_data = io_enq_bits_param;
  assign ram_param__T_29_addr = value;
  assign ram_param__T_29_mask = _T_25;
  assign ram_param__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_source__T_43_addr = value_1;
  assign ram_source__T_43_data = ram_source[ram_source__T_43_addr];
  assign ram_source__T_29_data = io_enq_bits_source;
  assign ram_source__T_29_addr = value;
  assign ram_source__T_29_mask = _T_25;
  assign ram_source__T_29_en = _T_25;
  assign ram_sink__T_43_addr = value_1;
  assign ram_sink__T_43_data = ram_sink[ram_sink__T_43_addr];
  assign ram_sink__T_29_data = io_enq_bits_sink;
  assign ram_sink__T_29_addr = value;
  assign ram_sink__T_29_mask = _T_25;
  assign ram_sink__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign ram_error__T_43_addr = value_1;
  assign ram_error__T_43_data = ram_error[ram_error__T_43_addr];
  assign ram_error__T_29_data = io_enq_bits_error;
  assign ram_error__T_29_addr = value;
  assign ram_error__T_29_mask = _T_25;
  assign ram_error__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_10 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_11 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_12 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_error[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_29_en & ram_opcode__T_29_mask) begin
      ram_opcode[ram_opcode__T_29_addr] <= ram_opcode__T_29_data;
    end
    if(ram_param__T_29_en & ram_param__T_29_mask) begin
      ram_param[ram_param__T_29_addr] <= ram_param__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_source__T_29_en & ram_source__T_29_mask) begin
      ram_source[ram_source__T_29_addr] <= ram_source__T_29_data;
    end
    if(ram_sink__T_29_en & ram_sink__T_29_mask) begin
      ram_sink[ram_sink__T_29_addr] <= ram_sink__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if(ram_error__T_29_en & ram_error__T_29_mask) begin
      ram_error[ram_error__T_29_addr] <= ram_error__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module TLBuffer_2(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [2:0] Queue_io_enq_bits_param;
  wire [2:0] Queue_io_enq_bits_size;
  wire [4:0] Queue_io_enq_bits_source;
  wire [31:0] Queue_io_enq_bits_address;
  wire [3:0] Queue_io_enq_bits_mask;
  wire [31:0] Queue_io_enq_bits_data;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [2:0] Queue_io_deq_bits_param;
  wire [2:0] Queue_io_deq_bits_size;
  wire [4:0] Queue_io_deq_bits_source;
  wire [31:0] Queue_io_deq_bits_address;
  wire [3:0] Queue_io_deq_bits_mask;
  wire [31:0] Queue_io_deq_bits_data;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [1:0] Queue_1_io_enq_bits_param;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [4:0] Queue_1_io_enq_bits_source;
  wire  Queue_1_io_enq_bits_sink;
  wire [31:0] Queue_1_io_enq_bits_data;
  wire  Queue_1_io_enq_bits_error;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [1:0] Queue_1_io_deq_bits_param;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [4:0] Queue_1_io_deq_bits_source;
  wire  Queue_1_io_deq_bits_sink;
  wire [31:0] Queue_1_io_deq_bits_data;
  wire  Queue_1_io_deq_bits_error;
  Queue_6 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_7 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_error(Queue_1_io_enq_bits_error),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_error(Queue_1_io_deq_bits_error)
  );
  assign io_in_0_a_ready = Queue_io_enq_ready;
  assign io_in_0_d_valid = Queue_1_io_deq_valid;
  assign io_in_0_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign io_in_0_d_bits_param = Queue_1_io_deq_bits_param;
  assign io_in_0_d_bits_size = Queue_1_io_deq_bits_size;
  assign io_in_0_d_bits_source = Queue_1_io_deq_bits_source;
  assign io_in_0_d_bits_sink = Queue_1_io_deq_bits_sink;
  assign io_in_0_d_bits_data = Queue_1_io_deq_bits_data;
  assign io_in_0_d_bits_error = Queue_1_io_deq_bits_error;
  assign io_out_0_a_valid = Queue_io_deq_valid;
  assign io_out_0_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign io_out_0_a_bits_param = Queue_io_deq_bits_param;
  assign io_out_0_a_bits_size = Queue_io_deq_bits_size;
  assign io_out_0_a_bits_source = Queue_io_deq_bits_source;
  assign io_out_0_a_bits_address = Queue_io_deq_bits_address;
  assign io_out_0_a_bits_mask = Queue_io_deq_bits_mask;
  assign io_out_0_a_bits_data = Queue_io_deq_bits_data;
  assign io_out_0_d_ready = Queue_1_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_a_valid;
  assign Queue_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Queue_io_enq_bits_param = io_in_0_a_bits_param;
  assign Queue_io_enq_bits_size = io_in_0_a_bits_size;
  assign Queue_io_enq_bits_source = io_in_0_a_bits_source;
  assign Queue_io_enq_bits_address = io_in_0_a_bits_address;
  assign Queue_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Queue_io_enq_bits_data = io_in_0_a_bits_data;
  assign Queue_io_deq_ready = io_out_0_a_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_out_0_d_valid;
  assign Queue_1_io_enq_bits_opcode = io_out_0_d_bits_opcode;
  assign Queue_1_io_enq_bits_param = io_out_0_d_bits_param;
  assign Queue_1_io_enq_bits_size = io_out_0_d_bits_size;
  assign Queue_1_io_enq_bits_source = io_out_0_d_bits_source;
  assign Queue_1_io_enq_bits_sink = io_out_0_d_bits_sink;
  assign Queue_1_io_enq_bits_data = io_out_0_d_bits_data;
  assign Queue_1_io_enq_bits_error = io_out_0_d_bits_error;
  assign Queue_1_io_deq_ready = io_in_0_d_ready;
endmodule
module TLBuffer_3(
  output        io_in_4_a_ready,
  input         io_in_4_a_valid,
  input  [2:0]  io_in_4_a_bits_opcode,
  input  [2:0]  io_in_4_a_bits_param,
  input  [2:0]  io_in_4_a_bits_size,
  input  [4:0]  io_in_4_a_bits_source,
  input  [31:0] io_in_4_a_bits_address,
  input  [3:0]  io_in_4_a_bits_mask,
  input  [31:0] io_in_4_a_bits_data,
  input         io_in_4_d_ready,
  output        io_in_4_d_valid,
  output [2:0]  io_in_4_d_bits_opcode,
  output [1:0]  io_in_4_d_bits_param,
  output [2:0]  io_in_4_d_bits_size,
  output [4:0]  io_in_4_d_bits_source,
  output        io_in_4_d_bits_sink,
  output [31:0] io_in_4_d_bits_data,
  output        io_in_4_d_bits_error,
  output        io_in_3_a_ready,
  input         io_in_3_a_valid,
  input  [2:0]  io_in_3_a_bits_opcode,
  input  [2:0]  io_in_3_a_bits_size,
  input  [4:0]  io_in_3_a_bits_source,
  input  [16:0] io_in_3_a_bits_address,
  input  [3:0]  io_in_3_a_bits_mask,
  input         io_in_3_d_ready,
  output        io_in_3_d_valid,
  output [2:0]  io_in_3_d_bits_opcode,
  output [1:0]  io_in_3_d_bits_param,
  output [2:0]  io_in_3_d_bits_size,
  output [4:0]  io_in_3_d_bits_source,
  output        io_in_3_d_bits_sink,
  output [31:0] io_in_3_d_bits_data,
  output        io_in_3_d_bits_error,
  output        io_in_2_a_ready,
  input         io_in_2_a_valid,
  input  [2:0]  io_in_2_a_bits_opcode,
  input  [2:0]  io_in_2_a_bits_size,
  input  [4:0]  io_in_2_a_bits_source,
  input  [11:0] io_in_2_a_bits_address,
  input  [3:0]  io_in_2_a_bits_mask,
  input  [31:0] io_in_2_a_bits_data,
  input         io_in_2_d_ready,
  output        io_in_2_d_valid,
  output [2:0]  io_in_2_d_bits_opcode,
  output [1:0]  io_in_2_d_bits_param,
  output [2:0]  io_in_2_d_bits_size,
  output [4:0]  io_in_2_d_bits_source,
  output        io_in_2_d_bits_sink,
  output [31:0] io_in_2_d_bits_data,
  output        io_in_2_d_bits_error,
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [2:0]  io_in_1_a_bits_size,
  input  [4:0]  io_in_1_a_bits_source,
  input  [25:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [1:0]  io_in_1_d_bits_param,
  output [2:0]  io_in_1_d_bits_size,
  output [4:0]  io_in_1_d_bits_source,
  output        io_in_1_d_bits_sink,
  output [31:0] io_in_1_d_bits_data,
  output        io_in_1_d_bits_error,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [27:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_4_a_ready,
  output        io_out_4_a_valid,
  output [2:0]  io_out_4_a_bits_opcode,
  output [2:0]  io_out_4_a_bits_param,
  output [2:0]  io_out_4_a_bits_size,
  output [4:0]  io_out_4_a_bits_source,
  output [31:0] io_out_4_a_bits_address,
  output [3:0]  io_out_4_a_bits_mask,
  output [31:0] io_out_4_a_bits_data,
  output        io_out_4_d_ready,
  input         io_out_4_d_valid,
  input  [2:0]  io_out_4_d_bits_opcode,
  input  [1:0]  io_out_4_d_bits_param,
  input  [2:0]  io_out_4_d_bits_size,
  input  [4:0]  io_out_4_d_bits_source,
  input         io_out_4_d_bits_sink,
  input  [31:0] io_out_4_d_bits_data,
  input         io_out_4_d_bits_error,
  input         io_out_3_a_ready,
  output        io_out_3_a_valid,
  output [2:0]  io_out_3_a_bits_opcode,
  output [2:0]  io_out_3_a_bits_size,
  output [4:0]  io_out_3_a_bits_source,
  output [16:0] io_out_3_a_bits_address,
  output [3:0]  io_out_3_a_bits_mask,
  output        io_out_3_d_ready,
  input         io_out_3_d_valid,
  input  [2:0]  io_out_3_d_bits_opcode,
  input  [1:0]  io_out_3_d_bits_param,
  input  [2:0]  io_out_3_d_bits_size,
  input  [4:0]  io_out_3_d_bits_source,
  input         io_out_3_d_bits_sink,
  input  [31:0] io_out_3_d_bits_data,
  input         io_out_3_d_bits_error,
  input         io_out_2_a_ready,
  output        io_out_2_a_valid,
  output [2:0]  io_out_2_a_bits_opcode,
  output [2:0]  io_out_2_a_bits_size,
  output [4:0]  io_out_2_a_bits_source,
  output [11:0] io_out_2_a_bits_address,
  output [3:0]  io_out_2_a_bits_mask,
  output [31:0] io_out_2_a_bits_data,
  output        io_out_2_d_ready,
  input         io_out_2_d_valid,
  input  [2:0]  io_out_2_d_bits_opcode,
  input  [1:0]  io_out_2_d_bits_param,
  input  [2:0]  io_out_2_d_bits_size,
  input  [4:0]  io_out_2_d_bits_source,
  input         io_out_2_d_bits_sink,
  input  [31:0] io_out_2_d_bits_data,
  input         io_out_2_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [2:0]  io_out_1_a_bits_size,
  output [4:0]  io_out_1_a_bits_source,
  output [25:0] io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [2:0]  io_out_1_d_bits_size,
  input  [4:0]  io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [31:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [27:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  assign io_in_4_a_ready = io_out_4_a_ready;
  assign io_in_4_d_valid = io_out_4_d_valid;
  assign io_in_4_d_bits_opcode = io_out_4_d_bits_opcode;
  assign io_in_4_d_bits_param = io_out_4_d_bits_param;
  assign io_in_4_d_bits_size = io_out_4_d_bits_size;
  assign io_in_4_d_bits_source = io_out_4_d_bits_source;
  assign io_in_4_d_bits_sink = io_out_4_d_bits_sink;
  assign io_in_4_d_bits_data = io_out_4_d_bits_data;
  assign io_in_4_d_bits_error = io_out_4_d_bits_error;
  assign io_in_3_a_ready = io_out_3_a_ready;
  assign io_in_3_d_valid = io_out_3_d_valid;
  assign io_in_3_d_bits_opcode = io_out_3_d_bits_opcode;
  assign io_in_3_d_bits_param = io_out_3_d_bits_param;
  assign io_in_3_d_bits_size = io_out_3_d_bits_size;
  assign io_in_3_d_bits_source = io_out_3_d_bits_source;
  assign io_in_3_d_bits_sink = io_out_3_d_bits_sink;
  assign io_in_3_d_bits_data = io_out_3_d_bits_data;
  assign io_in_3_d_bits_error = io_out_3_d_bits_error;
  assign io_in_2_a_ready = io_out_2_a_ready;
  assign io_in_2_d_valid = io_out_2_d_valid;
  assign io_in_2_d_bits_opcode = io_out_2_d_bits_opcode;
  assign io_in_2_d_bits_param = io_out_2_d_bits_param;
  assign io_in_2_d_bits_size = io_out_2_d_bits_size;
  assign io_in_2_d_bits_source = io_out_2_d_bits_source;
  assign io_in_2_d_bits_sink = io_out_2_d_bits_sink;
  assign io_in_2_d_bits_data = io_out_2_d_bits_data;
  assign io_in_2_d_bits_error = io_out_2_d_bits_error;
  assign io_in_1_a_ready = io_out_1_a_ready;
  assign io_in_1_d_valid = io_out_1_d_valid;
  assign io_in_1_d_bits_opcode = io_out_1_d_bits_opcode;
  assign io_in_1_d_bits_param = io_out_1_d_bits_param;
  assign io_in_1_d_bits_size = io_out_1_d_bits_size;
  assign io_in_1_d_bits_source = io_out_1_d_bits_source;
  assign io_in_1_d_bits_sink = io_out_1_d_bits_sink;
  assign io_in_1_d_bits_data = io_out_1_d_bits_data;
  assign io_in_1_d_bits_error = io_out_1_d_bits_error;
  assign io_in_0_a_ready = io_out_0_a_ready;
  assign io_in_0_d_valid = io_out_0_d_valid;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_param = io_out_0_d_bits_param;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_in_0_d_bits_sink = io_out_0_d_bits_sink;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_d_bits_error = io_out_0_d_bits_error;
  assign io_out_4_a_valid = io_in_4_a_valid;
  assign io_out_4_a_bits_opcode = io_in_4_a_bits_opcode;
  assign io_out_4_a_bits_param = io_in_4_a_bits_param;
  assign io_out_4_a_bits_size = io_in_4_a_bits_size;
  assign io_out_4_a_bits_source = io_in_4_a_bits_source;
  assign io_out_4_a_bits_address = io_in_4_a_bits_address;
  assign io_out_4_a_bits_mask = io_in_4_a_bits_mask;
  assign io_out_4_a_bits_data = io_in_4_a_bits_data;
  assign io_out_4_d_ready = io_in_4_d_ready;
  assign io_out_3_a_valid = io_in_3_a_valid;
  assign io_out_3_a_bits_opcode = io_in_3_a_bits_opcode;
  assign io_out_3_a_bits_size = io_in_3_a_bits_size;
  assign io_out_3_a_bits_source = io_in_3_a_bits_source;
  assign io_out_3_a_bits_address = io_in_3_a_bits_address;
  assign io_out_3_a_bits_mask = io_in_3_a_bits_mask;
  assign io_out_3_d_ready = io_in_3_d_ready;
  assign io_out_2_a_valid = io_in_2_a_valid;
  assign io_out_2_a_bits_opcode = io_in_2_a_bits_opcode;
  assign io_out_2_a_bits_size = io_in_2_a_bits_size;
  assign io_out_2_a_bits_source = io_in_2_a_bits_source;
  assign io_out_2_a_bits_address = io_in_2_a_bits_address;
  assign io_out_2_a_bits_mask = io_in_2_a_bits_mask;
  assign io_out_2_a_bits_data = io_in_2_a_bits_data;
  assign io_out_2_d_ready = io_in_2_d_ready;
  assign io_out_1_a_valid = io_in_1_a_valid;
  assign io_out_1_a_bits_opcode = io_in_1_a_bits_opcode;
  assign io_out_1_a_bits_size = io_in_1_a_bits_size;
  assign io_out_1_a_bits_source = io_in_1_a_bits_source;
  assign io_out_1_a_bits_address = io_in_1_a_bits_address;
  assign io_out_1_a_bits_mask = io_in_1_a_bits_mask;
  assign io_out_1_a_bits_data = io_in_1_a_bits_data;
  assign io_out_1_d_ready = io_in_1_d_ready;
  assign io_out_0_a_valid = io_in_0_a_valid;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address;
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = io_in_0_d_ready;
endmodule
module Repeater_1(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [27:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [27:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] saved_size;
  reg [31:0] _RAND_2;
  reg [4:0] saved_source;
  reg [31:0] _RAND_3;
  reg [27:0] saved_address;
  reg [31:0] _RAND_4;
  reg [3:0] saved_mask;
  reg [31:0] _RAND_5;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [2:0] _T_20_size;
  wire [4:0] _T_20_source;
  wire [27:0] _T_20_address;
  wire [3:0] _T_20_mask;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire [27:0] _GEN_5;
  wire [3:0] _GEN_6;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_full = full;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_address = _T_20_address;
  assign io_deq_bits_mask = _T_20_mask;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_address = full ? saved_address : io_enq_bits_address;
  assign _T_20_mask = full ? saved_mask : io_enq_bits_mask;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_address : saved_address;
  assign _GEN_6 = _T_22 ? io_enq_bits_mask : saved_mask;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_size = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_source = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_address = _RAND_4[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_mask = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_22) begin
      saved_mask <= io_enq_bits_mask;
    end
  end
endmodule
module Repeater_2(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [25:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [25:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] saved_size;
  reg [31:0] _RAND_2;
  reg [4:0] saved_source;
  reg [31:0] _RAND_3;
  reg [25:0] saved_address;
  reg [31:0] _RAND_4;
  reg [3:0] saved_mask;
  reg [31:0] _RAND_5;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [2:0] _T_20_size;
  wire [4:0] _T_20_source;
  wire [25:0] _T_20_address;
  wire [3:0] _T_20_mask;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire [25:0] _GEN_5;
  wire [3:0] _GEN_6;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_full = full;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_address = _T_20_address;
  assign io_deq_bits_mask = _T_20_mask;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_address = full ? saved_address : io_enq_bits_address;
  assign _T_20_mask = full ? saved_mask : io_enq_bits_mask;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_address : saved_address;
  assign _GEN_6 = _T_22 ? io_enq_bits_mask : saved_mask;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_size = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_source = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_address = _RAND_4[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_mask = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_22) begin
      saved_mask <= io_enq_bits_mask;
    end
  end
endmodule
module Repeater_3(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [11:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [11:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] saved_size;
  reg [31:0] _RAND_2;
  reg [4:0] saved_source;
  reg [31:0] _RAND_3;
  reg [11:0] saved_address;
  reg [31:0] _RAND_4;
  reg [3:0] saved_mask;
  reg [31:0] _RAND_5;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [2:0] _T_20_size;
  wire [4:0] _T_20_source;
  wire [11:0] _T_20_address;
  wire [3:0] _T_20_mask;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire [11:0] _GEN_5;
  wire [3:0] _GEN_6;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_full = full;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_address = _T_20_address;
  assign io_deq_bits_mask = _T_20_mask;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_address = full ? saved_address : io_enq_bits_address;
  assign _T_20_mask = full ? saved_mask : io_enq_bits_mask;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_address : saved_address;
  assign _GEN_6 = _T_22 ? io_enq_bits_mask : saved_mask;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_size = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_source = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_address = _RAND_4[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_mask = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_22) begin
      saved_mask <= io_enq_bits_mask;
    end
  end
endmodule
module Repeater_4(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [16:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [16:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] saved_size;
  reg [31:0] _RAND_2;
  reg [4:0] saved_source;
  reg [31:0] _RAND_3;
  reg [16:0] saved_address;
  reg [31:0] _RAND_4;
  reg [3:0] saved_mask;
  reg [31:0] _RAND_5;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [2:0] _T_20_size;
  wire [4:0] _T_20_source;
  wire [16:0] _T_20_address;
  wire [3:0] _T_20_mask;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire [16:0] _GEN_5;
  wire [3:0] _GEN_6;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_full = full;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_address = _T_20_address;
  assign io_deq_bits_mask = _T_20_mask;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_address = full ? saved_address : io_enq_bits_address;
  assign _T_20_mask = full ? saved_mask : io_enq_bits_mask;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_address : saved_address;
  assign _GEN_6 = _T_22 ? io_enq_bits_mask : saved_mask;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_size = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_source = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_address = _RAND_4[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_mask = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_22) begin
      saved_mask <= io_enq_bits_mask;
    end
  end
endmodule
module TLFragmenter_1(
  input         clock,
  input         reset,
  output        io_in_3_a_ready,
  input         io_in_3_a_valid,
  input  [2:0]  io_in_3_a_bits_opcode,
  input  [2:0]  io_in_3_a_bits_size,
  input  [4:0]  io_in_3_a_bits_source,
  input  [16:0] io_in_3_a_bits_address,
  input  [3:0]  io_in_3_a_bits_mask,
  input         io_in_3_d_ready,
  output        io_in_3_d_valid,
  output [2:0]  io_in_3_d_bits_opcode,
  output [1:0]  io_in_3_d_bits_param,
  output [2:0]  io_in_3_d_bits_size,
  output [4:0]  io_in_3_d_bits_source,
  output        io_in_3_d_bits_sink,
  output [31:0] io_in_3_d_bits_data,
  output        io_in_3_d_bits_error,
  output        io_in_2_a_ready,
  input         io_in_2_a_valid,
  input  [2:0]  io_in_2_a_bits_opcode,
  input  [2:0]  io_in_2_a_bits_size,
  input  [4:0]  io_in_2_a_bits_source,
  input  [11:0] io_in_2_a_bits_address,
  input  [3:0]  io_in_2_a_bits_mask,
  input  [31:0] io_in_2_a_bits_data,
  input         io_in_2_d_ready,
  output        io_in_2_d_valid,
  output [2:0]  io_in_2_d_bits_opcode,
  output [1:0]  io_in_2_d_bits_param,
  output [2:0]  io_in_2_d_bits_size,
  output [4:0]  io_in_2_d_bits_source,
  output        io_in_2_d_bits_sink,
  output [31:0] io_in_2_d_bits_data,
  output        io_in_2_d_bits_error,
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [2:0]  io_in_1_a_bits_size,
  input  [4:0]  io_in_1_a_bits_source,
  input  [25:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [1:0]  io_in_1_d_bits_param,
  output [2:0]  io_in_1_d_bits_size,
  output [4:0]  io_in_1_d_bits_source,
  output        io_in_1_d_bits_sink,
  output [31:0] io_in_1_d_bits_data,
  output        io_in_1_d_bits_error,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [27:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_3_a_ready,
  output        io_out_3_a_valid,
  output [1:0]  io_out_3_a_bits_size,
  output [9:0]  io_out_3_a_bits_source,
  output [16:0] io_out_3_a_bits_address,
  output        io_out_3_d_ready,
  input         io_out_3_d_valid,
  input  [2:0]  io_out_3_d_bits_opcode,
  input  [1:0]  io_out_3_d_bits_param,
  input  [1:0]  io_out_3_d_bits_size,
  input  [9:0]  io_out_3_d_bits_source,
  input         io_out_3_d_bits_sink,
  input  [31:0] io_out_3_d_bits_data,
  input         io_out_3_d_bits_error,
  input         io_out_2_a_ready,
  output        io_out_2_a_valid,
  output [2:0]  io_out_2_a_bits_opcode,
  output [1:0]  io_out_2_a_bits_size,
  output [9:0]  io_out_2_a_bits_source,
  output [11:0] io_out_2_a_bits_address,
  output [3:0]  io_out_2_a_bits_mask,
  output [31:0] io_out_2_a_bits_data,
  output        io_out_2_d_ready,
  input         io_out_2_d_valid,
  input  [2:0]  io_out_2_d_bits_opcode,
  input  [1:0]  io_out_2_d_bits_param,
  input  [1:0]  io_out_2_d_bits_size,
  input  [9:0]  io_out_2_d_bits_source,
  input         io_out_2_d_bits_sink,
  input  [31:0] io_out_2_d_bits_data,
  input         io_out_2_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [1:0]  io_out_1_a_bits_size,
  output [9:0]  io_out_1_a_bits_source,
  output [25:0] io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [1:0]  io_out_1_d_bits_size,
  input  [9:0]  io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [31:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [1:0]  io_out_0_a_bits_size,
  output [9:0]  io_out_0_a_bits_source,
  output [27:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [1:0]  io_out_0_d_bits_size,
  input  [9:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  reg [3:0] _T_353;
  reg [31:0] _RAND_0;
  reg [2:0] _T_355;
  reg [31:0] _RAND_1;
  reg  _T_358;
  reg [31:0] _RAND_2;
  wire [3:0] _T_359;
  wire  _T_361;
  wire  _T_363;
  wire [3:0] _T_366;
  wire [2:0] _T_367;
  wire [4:0] _T_370;
  wire [1:0] _T_371;
  wire [1:0] _T_372;
  wire  _T_373;
  wire  _T_389;
  wire  _T_390;
  wire [5:0] _GEN_32;
  wire [5:0] _T_391;
  wire [5:0] _GEN_33;
  wire [5:0] _T_392;
  wire [6:0] _GEN_34;
  wire [6:0] _T_393;
  wire [6:0] _T_395;
  wire [6:0] _T_397;
  wire [6:0] _T_398;
  wire [6:0] _T_399;
  wire [2:0] _T_400;
  wire [3:0] _T_401;
  wire  _T_403;
  wire [3:0] _GEN_35;
  wire [3:0] _T_404;
  wire [1:0] _T_405;
  wire [1:0] _T_406;
  wire  _T_408;
  wire [1:0] _T_409;
  wire  _T_410;
  wire [1:0] _T_411;
  wire [2:0] _T_412;
  wire  _T_413;
  wire [3:0] _GEN_36;
  wire [4:0] _T_414;
  wire [4:0] _T_415;
  wire [3:0] _T_416;
  wire [3:0] _T_417;
  wire  _T_418;
  wire [2:0] _GEN_0;
  wire  _GEN_1;
  wire [3:0] _GEN_2;
  wire [2:0] _GEN_3;
  wire  _GEN_4;
  wire  _T_420;
  wire  _T_422;
  wire  _T_423;
  wire  _T_424;
  wire  _T_426;
  wire  _T_427;
  wire [4:0] _T_428;
  reg  _T_432;
  reg [31:0] _RAND_3;
  wire  _T_433;
  wire  _T_436;
  wire  _GEN_5;
  wire  Repeater_clock;
  wire  Repeater_reset;
  wire  Repeater_io_repeat;
  wire  Repeater_io_full;
  wire  Repeater_io_enq_ready;
  wire  Repeater_io_enq_valid;
  wire [2:0] Repeater_io_enq_bits_opcode;
  wire [2:0] Repeater_io_enq_bits_size;
  wire [4:0] Repeater_io_enq_bits_source;
  wire [27:0] Repeater_io_enq_bits_address;
  wire [3:0] Repeater_io_enq_bits_mask;
  wire  Repeater_io_deq_ready;
  wire  Repeater_io_deq_valid;
  wire [2:0] Repeater_io_deq_bits_opcode;
  wire [2:0] Repeater_io_deq_bits_size;
  wire [4:0] Repeater_io_deq_bits_source;
  wire [27:0] Repeater_io_deq_bits_address;
  wire [3:0] Repeater_io_deq_bits_mask;
  wire  _T_473;
  wire [2:0] _T_474;
  wire [12:0] _T_477;
  wire [5:0] _T_478;
  wire [5:0] _T_479;
  wire [8:0] _T_482;
  wire [1:0] _T_483;
  wire [1:0] _T_484;
  wire  _T_485;
  wire  _T_487;
  reg [3:0] _T_492;
  reg [31:0] _RAND_4;
  wire  _T_494;
  wire [3:0] _T_495;
  wire [4:0] _T_497;
  wire [4:0] _T_498;
  wire [3:0] _T_499;
  wire [3:0] _T_500;
  wire [3:0] _T_501;
  wire [3:0] _T_504;
  reg  _T_513;
  reg [31:0] _RAND_5;
  wire  _GEN_6;
  wire  _T_516;
  wire  _T_517;
  wire [3:0] _GEN_7;
  wire  _T_519;
  wire  _T_521;
  wire  _T_522;
  wire [5:0] _GEN_37;
  wire [5:0] _T_523;
  wire [5:0] _T_524;
  wire [5:0] _T_525;
  wire [5:0] _GEN_38;
  wire [5:0] _T_526;
  wire [5:0] _T_528;
  wire [5:0] _T_529;
  wire [27:0] _GEN_39;
  wire [27:0] _T_530;
  wire [5:0] _T_531;
  wire [9:0] _T_532;
  wire  _T_534;
  wire  _T_537;
  wire  _T_538;
  wire  _T_540;
  wire  _T_544;
  wire  _T_545;
  wire  _T_546;
  wire  _T_548;
  wire [3:0] _T_549;
  reg [3:0] _T_558;
  reg [31:0] _RAND_6;
  reg [2:0] _T_560;
  reg [31:0] _RAND_7;
  reg  _T_563;
  reg [31:0] _RAND_8;
  wire [3:0] _T_564;
  wire  _T_566;
  wire  _T_568;
  wire [3:0] _T_571;
  wire [2:0] _T_572;
  wire [4:0] _T_575;
  wire [1:0] _T_576;
  wire [1:0] _T_577;
  wire  _T_578;
  wire  _T_594;
  wire  _T_595;
  wire [5:0] _GEN_40;
  wire [5:0] _T_596;
  wire [5:0] _GEN_41;
  wire [5:0] _T_597;
  wire [6:0] _GEN_42;
  wire [6:0] _T_598;
  wire [6:0] _T_600;
  wire [6:0] _T_602;
  wire [6:0] _T_603;
  wire [6:0] _T_604;
  wire [2:0] _T_605;
  wire [3:0] _T_606;
  wire  _T_608;
  wire [3:0] _GEN_43;
  wire [3:0] _T_609;
  wire [1:0] _T_610;
  wire [1:0] _T_611;
  wire  _T_613;
  wire [1:0] _T_614;
  wire  _T_615;
  wire [1:0] _T_616;
  wire [2:0] _T_617;
  wire  _T_618;
  wire [3:0] _GEN_44;
  wire [4:0] _T_619;
  wire [4:0] _T_620;
  wire [3:0] _T_621;
  wire [3:0] _T_622;
  wire  _T_623;
  wire [2:0] _GEN_8;
  wire  _GEN_9;
  wire [3:0] _GEN_10;
  wire [2:0] _GEN_11;
  wire  _GEN_12;
  wire  _T_625;
  wire  _T_627;
  wire  _T_628;
  wire  _T_629;
  wire  _T_631;
  wire  _T_632;
  wire [4:0] _T_633;
  reg  _T_637;
  reg [31:0] _RAND_9;
  wire  _T_638;
  wire  _T_641;
  wire  _GEN_13;
  wire  Repeater_1_clock;
  wire  Repeater_1_reset;
  wire  Repeater_1_io_repeat;
  wire  Repeater_1_io_full;
  wire  Repeater_1_io_enq_ready;
  wire  Repeater_1_io_enq_valid;
  wire [2:0] Repeater_1_io_enq_bits_opcode;
  wire [2:0] Repeater_1_io_enq_bits_size;
  wire [4:0] Repeater_1_io_enq_bits_source;
  wire [25:0] Repeater_1_io_enq_bits_address;
  wire [3:0] Repeater_1_io_enq_bits_mask;
  wire  Repeater_1_io_deq_ready;
  wire  Repeater_1_io_deq_valid;
  wire [2:0] Repeater_1_io_deq_bits_opcode;
  wire [2:0] Repeater_1_io_deq_bits_size;
  wire [4:0] Repeater_1_io_deq_bits_source;
  wire [25:0] Repeater_1_io_deq_bits_address;
  wire [3:0] Repeater_1_io_deq_bits_mask;
  wire  _T_678;
  wire [2:0] _T_679;
  wire [12:0] _T_682;
  wire [5:0] _T_683;
  wire [5:0] _T_684;
  wire [8:0] _T_687;
  wire [1:0] _T_688;
  wire [1:0] _T_689;
  wire  _T_690;
  wire  _T_692;
  reg [3:0] _T_697;
  reg [31:0] _RAND_10;
  wire  _T_699;
  wire [3:0] _T_700;
  wire [4:0] _T_702;
  wire [4:0] _T_703;
  wire [3:0] _T_704;
  wire [3:0] _T_705;
  wire [3:0] _T_706;
  wire [3:0] _T_709;
  reg  _T_718;
  reg [31:0] _RAND_11;
  wire  _GEN_14;
  wire  _T_721;
  wire  _T_722;
  wire [3:0] _GEN_15;
  wire  _T_724;
  wire  _T_726;
  wire  _T_727;
  wire [5:0] _GEN_45;
  wire [5:0] _T_728;
  wire [5:0] _T_729;
  wire [5:0] _T_730;
  wire [5:0] _GEN_46;
  wire [5:0] _T_731;
  wire [5:0] _T_733;
  wire [5:0] _T_734;
  wire [25:0] _GEN_47;
  wire [25:0] _T_735;
  wire [5:0] _T_736;
  wire [9:0] _T_737;
  wire  _T_739;
  wire  _T_742;
  wire  _T_743;
  wire  _T_745;
  wire  _T_749;
  wire  _T_750;
  wire  _T_751;
  wire  _T_753;
  wire [3:0] _T_754;
  reg [3:0] _T_763;
  reg [31:0] _RAND_12;
  reg [2:0] _T_765;
  reg [31:0] _RAND_13;
  reg  _T_768;
  reg [31:0] _RAND_14;
  wire [3:0] _T_769;
  wire  _T_771;
  wire  _T_773;
  wire [3:0] _T_776;
  wire [2:0] _T_777;
  wire [4:0] _T_780;
  wire [1:0] _T_781;
  wire [1:0] _T_782;
  wire  _T_783;
  wire  _T_799;
  wire  _T_800;
  wire [5:0] _GEN_48;
  wire [5:0] _T_801;
  wire [5:0] _GEN_49;
  wire [5:0] _T_802;
  wire [6:0] _GEN_50;
  wire [6:0] _T_803;
  wire [6:0] _T_805;
  wire [6:0] _T_807;
  wire [6:0] _T_808;
  wire [6:0] _T_809;
  wire [2:0] _T_810;
  wire [3:0] _T_811;
  wire  _T_813;
  wire [3:0] _GEN_51;
  wire [3:0] _T_814;
  wire [1:0] _T_815;
  wire [1:0] _T_816;
  wire  _T_818;
  wire [1:0] _T_819;
  wire  _T_820;
  wire [1:0] _T_821;
  wire [2:0] _T_822;
  wire  _T_823;
  wire [3:0] _GEN_52;
  wire [4:0] _T_824;
  wire [4:0] _T_825;
  wire [3:0] _T_826;
  wire [3:0] _T_827;
  wire  _T_828;
  wire [2:0] _GEN_16;
  wire  _GEN_17;
  wire [3:0] _GEN_18;
  wire [2:0] _GEN_19;
  wire  _GEN_20;
  wire  _T_830;
  wire  _T_832;
  wire  _T_833;
  wire  _T_834;
  wire  _T_836;
  wire  _T_837;
  wire [4:0] _T_838;
  reg  _T_842;
  reg [31:0] _RAND_15;
  wire  _T_843;
  wire  _T_846;
  wire  _GEN_21;
  wire  Repeater_2_clock;
  wire  Repeater_2_reset;
  wire  Repeater_2_io_repeat;
  wire  Repeater_2_io_full;
  wire  Repeater_2_io_enq_ready;
  wire  Repeater_2_io_enq_valid;
  wire [2:0] Repeater_2_io_enq_bits_opcode;
  wire [2:0] Repeater_2_io_enq_bits_size;
  wire [4:0] Repeater_2_io_enq_bits_source;
  wire [11:0] Repeater_2_io_enq_bits_address;
  wire [3:0] Repeater_2_io_enq_bits_mask;
  wire  Repeater_2_io_deq_ready;
  wire  Repeater_2_io_deq_valid;
  wire [2:0] Repeater_2_io_deq_bits_opcode;
  wire [2:0] Repeater_2_io_deq_bits_size;
  wire [4:0] Repeater_2_io_deq_bits_source;
  wire [11:0] Repeater_2_io_deq_bits_address;
  wire [3:0] Repeater_2_io_deq_bits_mask;
  wire  _T_883;
  wire [2:0] _T_884;
  wire [12:0] _T_887;
  wire [5:0] _T_888;
  wire [5:0] _T_889;
  wire [8:0] _T_892;
  wire [1:0] _T_893;
  wire [1:0] _T_894;
  wire  _T_895;
  wire  _T_897;
  reg [3:0] _T_902;
  reg [31:0] _RAND_16;
  wire  _T_904;
  wire [3:0] _T_905;
  wire [4:0] _T_907;
  wire [4:0] _T_908;
  wire [3:0] _T_909;
  wire [3:0] _T_910;
  wire [3:0] _T_911;
  wire [3:0] _T_914;
  reg  _T_923;
  reg [31:0] _RAND_17;
  wire  _GEN_22;
  wire  _T_926;
  wire  _T_927;
  wire [3:0] _GEN_23;
  wire  _T_929;
  wire  _T_931;
  wire  _T_932;
  wire [5:0] _GEN_53;
  wire [5:0] _T_933;
  wire [5:0] _T_934;
  wire [5:0] _T_935;
  wire [5:0] _GEN_54;
  wire [5:0] _T_936;
  wire [5:0] _T_938;
  wire [5:0] _T_939;
  wire [11:0] _GEN_55;
  wire [11:0] _T_940;
  wire [5:0] _T_941;
  wire [9:0] _T_942;
  wire  _T_944;
  wire  _T_947;
  wire  _T_948;
  wire  _T_950;
  wire  _T_954;
  wire  _T_955;
  wire  _T_956;
  wire  _T_958;
  wire [3:0] _T_959;
  reg [3:0] _T_968;
  reg [31:0] _RAND_18;
  reg [2:0] _T_970;
  reg [31:0] _RAND_19;
  reg  _T_973;
  reg [31:0] _RAND_20;
  wire [3:0] _T_974;
  wire  _T_976;
  wire [4:0] _T_985;
  wire [1:0] _T_986;
  wire [1:0] _T_987;
  wire [5:0] _GEN_56;
  wire [5:0] _T_1007;
  wire [5:0] _GEN_57;
  wire [5:0] _T_1008;
  wire [6:0] _GEN_58;
  wire [6:0] _T_1009;
  wire [6:0] _T_1011;
  wire [6:0] _T_1013;
  wire [6:0] _T_1014;
  wire [6:0] _T_1015;
  wire [2:0] _T_1016;
  wire [3:0] _T_1017;
  wire  _T_1019;
  wire [3:0] _GEN_59;
  wire [3:0] _T_1020;
  wire [1:0] _T_1021;
  wire [1:0] _T_1022;
  wire  _T_1024;
  wire [1:0] _T_1025;
  wire  _T_1026;
  wire [1:0] _T_1027;
  wire [2:0] _T_1028;
  wire  _T_1029;
  wire [4:0] _T_1030;
  wire [4:0] _T_1031;
  wire [3:0] _T_1032;
  wire [3:0] _T_1033;
  wire  _T_1034;
  wire [2:0] _GEN_24;
  wire  _GEN_25;
  wire [3:0] _GEN_26;
  wire [2:0] _GEN_27;
  wire  _GEN_28;
  wire [4:0] _T_1044;
  reg  _T_1048;
  reg [31:0] _RAND_21;
  wire  _T_1049;
  wire  _GEN_29;
  wire  Repeater_3_clock;
  wire  Repeater_3_reset;
  wire  Repeater_3_io_repeat;
  wire  Repeater_3_io_full;
  wire  Repeater_3_io_enq_ready;
  wire  Repeater_3_io_enq_valid;
  wire [2:0] Repeater_3_io_enq_bits_opcode;
  wire [2:0] Repeater_3_io_enq_bits_size;
  wire [4:0] Repeater_3_io_enq_bits_source;
  wire [16:0] Repeater_3_io_enq_bits_address;
  wire [3:0] Repeater_3_io_enq_bits_mask;
  wire  Repeater_3_io_deq_ready;
  wire  Repeater_3_io_deq_valid;
  wire [2:0] Repeater_3_io_deq_bits_opcode;
  wire [2:0] Repeater_3_io_deq_bits_size;
  wire [4:0] Repeater_3_io_deq_bits_source;
  wire [16:0] Repeater_3_io_deq_bits_address;
  wire [3:0] Repeater_3_io_deq_bits_mask;
  wire  _T_1087;
  wire [2:0] _T_1088;
  wire [12:0] _T_1091;
  wire [5:0] _T_1092;
  wire [5:0] _T_1093;
  wire [8:0] _T_1096;
  wire [1:0] _T_1097;
  wire [1:0] _T_1098;
  wire  _T_1099;
  wire  _T_1101;
  reg [3:0] _T_1106;
  reg [31:0] _RAND_22;
  wire  _T_1108;
  wire [3:0] _T_1109;
  wire [4:0] _T_1111;
  wire [4:0] _T_1112;
  wire [3:0] _T_1113;
  wire [3:0] _T_1114;
  wire [3:0] _T_1115;
  wire [3:0] _T_1118;
  reg  _T_1127;
  reg [31:0] _RAND_23;
  wire  _GEN_30;
  wire  _T_1130;
  wire  _T_1131;
  wire [3:0] _GEN_31;
  wire  _T_1133;
  wire  _T_1135;
  wire  _T_1136;
  wire [5:0] _GEN_60;
  wire [5:0] _T_1137;
  wire [5:0] _T_1138;
  wire [5:0] _T_1139;
  wire [5:0] _GEN_61;
  wire [5:0] _T_1140;
  wire [5:0] _T_1142;
  wire [5:0] _T_1143;
  wire [16:0] _GEN_62;
  wire [16:0] _T_1144;
  wire [5:0] _T_1145;
  wire [9:0] _T_1146;
  wire  _T_1148;
  wire  _T_1151;
  wire  _T_1152;
  wire  _T_1154;
  wire  _T_1158;
  wire  _T_1159;
  wire  _T_1160;
  wire  _T_1162;
  Repeater_1 Repeater (
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_full(Repeater_io_full),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_address(Repeater_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_io_enq_bits_mask),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_address(Repeater_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_io_deq_bits_mask)
  );
  Repeater_2 Repeater_1 (
    .clock(Repeater_1_clock),
    .reset(Repeater_1_reset),
    .io_repeat(Repeater_1_io_repeat),
    .io_full(Repeater_1_io_full),
    .io_enq_ready(Repeater_1_io_enq_ready),
    .io_enq_valid(Repeater_1_io_enq_valid),
    .io_enq_bits_opcode(Repeater_1_io_enq_bits_opcode),
    .io_enq_bits_size(Repeater_1_io_enq_bits_size),
    .io_enq_bits_source(Repeater_1_io_enq_bits_source),
    .io_enq_bits_address(Repeater_1_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_1_io_enq_bits_mask),
    .io_deq_ready(Repeater_1_io_deq_ready),
    .io_deq_valid(Repeater_1_io_deq_valid),
    .io_deq_bits_opcode(Repeater_1_io_deq_bits_opcode),
    .io_deq_bits_size(Repeater_1_io_deq_bits_size),
    .io_deq_bits_source(Repeater_1_io_deq_bits_source),
    .io_deq_bits_address(Repeater_1_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_1_io_deq_bits_mask)
  );
  Repeater_3 Repeater_2 (
    .clock(Repeater_2_clock),
    .reset(Repeater_2_reset),
    .io_repeat(Repeater_2_io_repeat),
    .io_full(Repeater_2_io_full),
    .io_enq_ready(Repeater_2_io_enq_ready),
    .io_enq_valid(Repeater_2_io_enq_valid),
    .io_enq_bits_opcode(Repeater_2_io_enq_bits_opcode),
    .io_enq_bits_size(Repeater_2_io_enq_bits_size),
    .io_enq_bits_source(Repeater_2_io_enq_bits_source),
    .io_enq_bits_address(Repeater_2_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_2_io_enq_bits_mask),
    .io_deq_ready(Repeater_2_io_deq_ready),
    .io_deq_valid(Repeater_2_io_deq_valid),
    .io_deq_bits_opcode(Repeater_2_io_deq_bits_opcode),
    .io_deq_bits_size(Repeater_2_io_deq_bits_size),
    .io_deq_bits_source(Repeater_2_io_deq_bits_source),
    .io_deq_bits_address(Repeater_2_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_2_io_deq_bits_mask)
  );
  Repeater_4 Repeater_3 (
    .clock(Repeater_3_clock),
    .reset(Repeater_3_reset),
    .io_repeat(Repeater_3_io_repeat),
    .io_full(Repeater_3_io_full),
    .io_enq_ready(Repeater_3_io_enq_ready),
    .io_enq_valid(Repeater_3_io_enq_valid),
    .io_enq_bits_opcode(Repeater_3_io_enq_bits_opcode),
    .io_enq_bits_size(Repeater_3_io_enq_bits_size),
    .io_enq_bits_source(Repeater_3_io_enq_bits_source),
    .io_enq_bits_address(Repeater_3_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_3_io_enq_bits_mask),
    .io_deq_ready(Repeater_3_io_deq_ready),
    .io_deq_valid(Repeater_3_io_deq_valid),
    .io_deq_bits_opcode(Repeater_3_io_deq_bits_opcode),
    .io_deq_bits_size(Repeater_3_io_deq_bits_size),
    .io_deq_bits_source(Repeater_3_io_deq_bits_source),
    .io_deq_bits_address(Repeater_3_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_3_io_deq_bits_mask)
  );
  assign io_in_3_a_ready = Repeater_3_io_enq_ready;
  assign io_in_3_d_valid = io_out_3_d_valid;
  assign io_in_3_d_bits_opcode = io_out_3_d_bits_opcode;
  assign io_in_3_d_bits_param = io_out_3_d_bits_param;
  assign io_in_3_d_bits_size = _GEN_24;
  assign io_in_3_d_bits_source = _T_1044;
  assign io_in_3_d_bits_sink = io_out_3_d_bits_sink;
  assign io_in_3_d_bits_data = io_out_3_d_bits_data;
  assign io_in_3_d_bits_error = _T_1049;
  assign io_in_2_a_ready = Repeater_2_io_enq_ready;
  assign io_in_2_d_valid = _T_837;
  assign io_in_2_d_bits_opcode = io_out_2_d_bits_opcode;
  assign io_in_2_d_bits_param = io_out_2_d_bits_param;
  assign io_in_2_d_bits_size = _GEN_16;
  assign io_in_2_d_bits_source = _T_838;
  assign io_in_2_d_bits_sink = io_out_2_d_bits_sink;
  assign io_in_2_d_bits_data = io_out_2_d_bits_data;
  assign io_in_2_d_bits_error = _T_843;
  assign io_in_1_a_ready = Repeater_1_io_enq_ready;
  assign io_in_1_d_valid = _T_632;
  assign io_in_1_d_bits_opcode = io_out_1_d_bits_opcode;
  assign io_in_1_d_bits_param = io_out_1_d_bits_param;
  assign io_in_1_d_bits_size = _GEN_8;
  assign io_in_1_d_bits_source = _T_633;
  assign io_in_1_d_bits_sink = io_out_1_d_bits_sink;
  assign io_in_1_d_bits_data = io_out_1_d_bits_data;
  assign io_in_1_d_bits_error = _T_638;
  assign io_in_0_a_ready = Repeater_io_enq_ready;
  assign io_in_0_d_valid = _T_427;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_param = io_out_0_d_bits_param;
  assign io_in_0_d_bits_size = _GEN_0;
  assign io_in_0_d_bits_source = _T_428;
  assign io_in_0_d_bits_sink = io_out_0_d_bits_sink;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_d_bits_error = _T_433;
  assign io_out_3_a_valid = Repeater_3_io_deq_valid;
  assign io_out_3_a_bits_size = _T_1088[1:0];
  assign io_out_3_a_bits_source = _T_1146;
  assign io_out_3_a_bits_address = _T_1144;
  assign io_out_3_d_ready = io_in_3_d_ready;
  assign io_out_2_a_valid = Repeater_2_io_deq_valid;
  assign io_out_2_a_bits_opcode = Repeater_2_io_deq_bits_opcode;
  assign io_out_2_a_bits_size = _T_884[1:0];
  assign io_out_2_a_bits_source = _T_942;
  assign io_out_2_a_bits_address = _T_940;
  assign io_out_2_a_bits_mask = _T_959;
  assign io_out_2_a_bits_data = io_in_2_a_bits_data;
  assign io_out_2_d_ready = _T_834;
  assign io_out_1_a_valid = Repeater_1_io_deq_valid;
  assign io_out_1_a_bits_opcode = Repeater_1_io_deq_bits_opcode;
  assign io_out_1_a_bits_size = _T_679[1:0];
  assign io_out_1_a_bits_source = _T_737;
  assign io_out_1_a_bits_address = _T_735;
  assign io_out_1_a_bits_mask = _T_754;
  assign io_out_1_a_bits_data = io_in_1_a_bits_data;
  assign io_out_1_d_ready = _T_629;
  assign io_out_0_a_valid = Repeater_io_deq_valid;
  assign io_out_0_a_bits_opcode = Repeater_io_deq_bits_opcode;
  assign io_out_0_a_bits_size = _T_474[1:0];
  assign io_out_0_a_bits_source = _T_532;
  assign io_out_0_a_bits_address = _T_530;
  assign io_out_0_a_bits_mask = _T_549;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = _T_424;
  assign _T_359 = io_out_0_d_bits_source[3:0];
  assign _T_361 = _T_353 == 4'h0;
  assign _T_363 = _T_359 == 4'h0;
  assign _T_366 = 4'h1 << io_out_0_d_bits_size;
  assign _T_367 = _T_366[2:0];
  assign _T_370 = 5'h3 << io_out_0_d_bits_size;
  assign _T_371 = _T_370[1:0];
  assign _T_372 = ~ _T_371;
  assign _T_373 = io_out_0_d_bits_opcode[0];
  assign _T_389 = _T_367[2:2];
  assign _T_390 = _T_373 ? 1'h1 : _T_389;
  assign _GEN_32 = {{2'd0}, _T_359};
  assign _T_391 = _GEN_32 << 2;
  assign _GEN_33 = {{4'd0}, _T_372};
  assign _T_392 = _T_391 | _GEN_33;
  assign _GEN_34 = {{1'd0}, _T_392};
  assign _T_393 = _GEN_34 << 1;
  assign _T_395 = _T_393 | 7'h1;
  assign _T_397 = {1'h0,_T_392};
  assign _T_398 = ~ _T_397;
  assign _T_399 = _T_395 & _T_398;
  assign _T_400 = _T_399[6:4];
  assign _T_401 = _T_399[3:0];
  assign _T_403 = _T_400 != 3'h0;
  assign _GEN_35 = {{1'd0}, _T_400};
  assign _T_404 = _GEN_35 | _T_401;
  assign _T_405 = _T_404[3:2];
  assign _T_406 = _T_404[1:0];
  assign _T_408 = _T_405 != 2'h0;
  assign _T_409 = _T_405 | _T_406;
  assign _T_410 = _T_409[1];
  assign _T_411 = {_T_408,_T_410};
  assign _T_412 = {_T_403,_T_411};
  assign _T_413 = io_out_0_d_ready & io_out_0_d_valid;
  assign _GEN_36 = {{3'd0}, _T_390};
  assign _T_414 = _T_353 - _GEN_36;
  assign _T_415 = $unsigned(_T_414);
  assign _T_416 = _T_415[3:0];
  assign _T_417 = _T_361 ? _T_359 : _T_416;
  assign _T_418 = io_out_0_d_bits_source[4];
  assign _GEN_0 = _T_361 ? _T_412 : _T_355;
  assign _GEN_1 = _T_361 ? _T_418 : _T_358;
  assign _GEN_2 = _T_413 ? _T_417 : _T_353;
  assign _GEN_3 = _T_413 ? _GEN_0 : _T_355;
  assign _GEN_4 = _T_413 ? _GEN_1 : _T_358;
  assign _T_420 = _T_373 == 1'h0;
  assign _T_422 = _T_363 == 1'h0;
  assign _T_423 = _T_420 & _T_422;
  assign _T_424 = io_in_0_d_ready | _T_423;
  assign _T_426 = _T_423 == 1'h0;
  assign _T_427 = io_out_0_d_valid & _T_426;
  assign _T_428 = io_out_0_d_bits_source[9:5];
  assign _T_433 = _T_432 | io_out_0_d_bits_error;
  assign _T_436 = _T_423 ? _T_433 : 1'h0;
  assign _GEN_5 = _T_413 ? _T_436 : _T_432;
  assign Repeater_clock = clock;
  assign Repeater_reset = reset;
  assign Repeater_io_repeat = _T_522;
  assign Repeater_io_enq_valid = io_in_0_a_valid;
  assign Repeater_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Repeater_io_enq_bits_size = io_in_0_a_bits_size;
  assign Repeater_io_enq_bits_source = io_in_0_a_bits_source;
  assign Repeater_io_enq_bits_address = io_in_0_a_bits_address;
  assign Repeater_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Repeater_io_deq_ready = io_out_0_a_ready;
  assign _T_473 = Repeater_io_deq_bits_size > 3'h2;
  assign _T_474 = _T_473 ? 3'h2 : Repeater_io_deq_bits_size;
  assign _T_477 = 13'h3f << Repeater_io_deq_bits_size;
  assign _T_478 = _T_477[5:0];
  assign _T_479 = ~ _T_478;
  assign _T_482 = 9'h3 << _T_474;
  assign _T_483 = _T_482[1:0];
  assign _T_484 = ~ _T_483;
  assign _T_485 = Repeater_io_deq_bits_opcode[2];
  assign _T_487 = _T_485 == 1'h0;
  assign _T_494 = _T_492 == 4'h0;
  assign _T_495 = _T_479[5:2];
  assign _T_497 = _T_492 - 4'h1;
  assign _T_498 = $unsigned(_T_497);
  assign _T_499 = _T_498[3:0];
  assign _T_500 = _T_494 ? _T_495 : _T_499;
  assign _T_501 = ~ _T_500;
  assign _T_504 = ~ _T_501;
  assign _GEN_6 = _T_494 ? _T_358 : _T_513;
  assign _T_516 = _GEN_6 == 1'h0;
  assign _T_517 = io_out_0_a_ready & io_out_0_a_valid;
  assign _GEN_7 = _T_517 ? _T_504 : _T_492;
  assign _T_519 = _T_487 == 1'h0;
  assign _T_521 = _T_504 != 4'h0;
  assign _T_522 = _T_519 & _T_521;
  assign _GEN_37 = {{2'd0}, _T_500};
  assign _T_523 = _GEN_37 << 2;
  assign _T_524 = ~ _T_479;
  assign _T_525 = _T_523 | _T_524;
  assign _GEN_38 = {{4'd0}, _T_484};
  assign _T_526 = _T_525 | _GEN_38;
  assign _T_528 = _T_526 | 6'h3;
  assign _T_529 = ~ _T_528;
  assign _GEN_39 = {{22'd0}, _T_529};
  assign _T_530 = Repeater_io_deq_bits_address | _GEN_39;
  assign _T_531 = {Repeater_io_deq_bits_source,_T_516};
  assign _T_532 = {_T_531,_T_504};
  assign _T_534 = Repeater_io_full == 1'h0;
  assign _T_537 = _T_534 | _T_519;
  assign _T_538 = _T_537 | reset;
  assign _T_540 = _T_538 == 1'h0;
  assign _T_544 = Repeater_io_deq_bits_mask == 4'hf;
  assign _T_545 = _T_534 | _T_544;
  assign _T_546 = _T_545 | reset;
  assign _T_548 = _T_546 == 1'h0;
  assign _T_549 = Repeater_io_full ? 4'hf : io_in_0_a_bits_mask;
  assign _T_564 = io_out_1_d_bits_source[3:0];
  assign _T_566 = _T_558 == 4'h0;
  assign _T_568 = _T_564 == 4'h0;
  assign _T_571 = 4'h1 << io_out_1_d_bits_size;
  assign _T_572 = _T_571[2:0];
  assign _T_575 = 5'h3 << io_out_1_d_bits_size;
  assign _T_576 = _T_575[1:0];
  assign _T_577 = ~ _T_576;
  assign _T_578 = io_out_1_d_bits_opcode[0];
  assign _T_594 = _T_572[2:2];
  assign _T_595 = _T_578 ? 1'h1 : _T_594;
  assign _GEN_40 = {{2'd0}, _T_564};
  assign _T_596 = _GEN_40 << 2;
  assign _GEN_41 = {{4'd0}, _T_577};
  assign _T_597 = _T_596 | _GEN_41;
  assign _GEN_42 = {{1'd0}, _T_597};
  assign _T_598 = _GEN_42 << 1;
  assign _T_600 = _T_598 | 7'h1;
  assign _T_602 = {1'h0,_T_597};
  assign _T_603 = ~ _T_602;
  assign _T_604 = _T_600 & _T_603;
  assign _T_605 = _T_604[6:4];
  assign _T_606 = _T_604[3:0];
  assign _T_608 = _T_605 != 3'h0;
  assign _GEN_43 = {{1'd0}, _T_605};
  assign _T_609 = _GEN_43 | _T_606;
  assign _T_610 = _T_609[3:2];
  assign _T_611 = _T_609[1:0];
  assign _T_613 = _T_610 != 2'h0;
  assign _T_614 = _T_610 | _T_611;
  assign _T_615 = _T_614[1];
  assign _T_616 = {_T_613,_T_615};
  assign _T_617 = {_T_608,_T_616};
  assign _T_618 = io_out_1_d_ready & io_out_1_d_valid;
  assign _GEN_44 = {{3'd0}, _T_595};
  assign _T_619 = _T_558 - _GEN_44;
  assign _T_620 = $unsigned(_T_619);
  assign _T_621 = _T_620[3:0];
  assign _T_622 = _T_566 ? _T_564 : _T_621;
  assign _T_623 = io_out_1_d_bits_source[4];
  assign _GEN_8 = _T_566 ? _T_617 : _T_560;
  assign _GEN_9 = _T_566 ? _T_623 : _T_563;
  assign _GEN_10 = _T_618 ? _T_622 : _T_558;
  assign _GEN_11 = _T_618 ? _GEN_8 : _T_560;
  assign _GEN_12 = _T_618 ? _GEN_9 : _T_563;
  assign _T_625 = _T_578 == 1'h0;
  assign _T_627 = _T_568 == 1'h0;
  assign _T_628 = _T_625 & _T_627;
  assign _T_629 = io_in_1_d_ready | _T_628;
  assign _T_631 = _T_628 == 1'h0;
  assign _T_632 = io_out_1_d_valid & _T_631;
  assign _T_633 = io_out_1_d_bits_source[9:5];
  assign _T_638 = _T_637 | io_out_1_d_bits_error;
  assign _T_641 = _T_628 ? _T_638 : 1'h0;
  assign _GEN_13 = _T_618 ? _T_641 : _T_637;
  assign Repeater_1_clock = clock;
  assign Repeater_1_reset = reset;
  assign Repeater_1_io_repeat = _T_727;
  assign Repeater_1_io_enq_valid = io_in_1_a_valid;
  assign Repeater_1_io_enq_bits_opcode = io_in_1_a_bits_opcode;
  assign Repeater_1_io_enq_bits_size = io_in_1_a_bits_size;
  assign Repeater_1_io_enq_bits_source = io_in_1_a_bits_source;
  assign Repeater_1_io_enq_bits_address = io_in_1_a_bits_address;
  assign Repeater_1_io_enq_bits_mask = io_in_1_a_bits_mask;
  assign Repeater_1_io_deq_ready = io_out_1_a_ready;
  assign _T_678 = Repeater_1_io_deq_bits_size > 3'h2;
  assign _T_679 = _T_678 ? 3'h2 : Repeater_1_io_deq_bits_size;
  assign _T_682 = 13'h3f << Repeater_1_io_deq_bits_size;
  assign _T_683 = _T_682[5:0];
  assign _T_684 = ~ _T_683;
  assign _T_687 = 9'h3 << _T_679;
  assign _T_688 = _T_687[1:0];
  assign _T_689 = ~ _T_688;
  assign _T_690 = Repeater_1_io_deq_bits_opcode[2];
  assign _T_692 = _T_690 == 1'h0;
  assign _T_699 = _T_697 == 4'h0;
  assign _T_700 = _T_684[5:2];
  assign _T_702 = _T_697 - 4'h1;
  assign _T_703 = $unsigned(_T_702);
  assign _T_704 = _T_703[3:0];
  assign _T_705 = _T_699 ? _T_700 : _T_704;
  assign _T_706 = ~ _T_705;
  assign _T_709 = ~ _T_706;
  assign _GEN_14 = _T_699 ? _T_563 : _T_718;
  assign _T_721 = _GEN_14 == 1'h0;
  assign _T_722 = io_out_1_a_ready & io_out_1_a_valid;
  assign _GEN_15 = _T_722 ? _T_709 : _T_697;
  assign _T_724 = _T_692 == 1'h0;
  assign _T_726 = _T_709 != 4'h0;
  assign _T_727 = _T_724 & _T_726;
  assign _GEN_45 = {{2'd0}, _T_705};
  assign _T_728 = _GEN_45 << 2;
  assign _T_729 = ~ _T_684;
  assign _T_730 = _T_728 | _T_729;
  assign _GEN_46 = {{4'd0}, _T_689};
  assign _T_731 = _T_730 | _GEN_46;
  assign _T_733 = _T_731 | 6'h3;
  assign _T_734 = ~ _T_733;
  assign _GEN_47 = {{20'd0}, _T_734};
  assign _T_735 = Repeater_1_io_deq_bits_address | _GEN_47;
  assign _T_736 = {Repeater_1_io_deq_bits_source,_T_721};
  assign _T_737 = {_T_736,_T_709};
  assign _T_739 = Repeater_1_io_full == 1'h0;
  assign _T_742 = _T_739 | _T_724;
  assign _T_743 = _T_742 | reset;
  assign _T_745 = _T_743 == 1'h0;
  assign _T_749 = Repeater_1_io_deq_bits_mask == 4'hf;
  assign _T_750 = _T_739 | _T_749;
  assign _T_751 = _T_750 | reset;
  assign _T_753 = _T_751 == 1'h0;
  assign _T_754 = Repeater_1_io_full ? 4'hf : io_in_1_a_bits_mask;
  assign _T_769 = io_out_2_d_bits_source[3:0];
  assign _T_771 = _T_763 == 4'h0;
  assign _T_773 = _T_769 == 4'h0;
  assign _T_776 = 4'h1 << io_out_2_d_bits_size;
  assign _T_777 = _T_776[2:0];
  assign _T_780 = 5'h3 << io_out_2_d_bits_size;
  assign _T_781 = _T_780[1:0];
  assign _T_782 = ~ _T_781;
  assign _T_783 = io_out_2_d_bits_opcode[0];
  assign _T_799 = _T_777[2:2];
  assign _T_800 = _T_783 ? 1'h1 : _T_799;
  assign _GEN_48 = {{2'd0}, _T_769};
  assign _T_801 = _GEN_48 << 2;
  assign _GEN_49 = {{4'd0}, _T_782};
  assign _T_802 = _T_801 | _GEN_49;
  assign _GEN_50 = {{1'd0}, _T_802};
  assign _T_803 = _GEN_50 << 1;
  assign _T_805 = _T_803 | 7'h1;
  assign _T_807 = {1'h0,_T_802};
  assign _T_808 = ~ _T_807;
  assign _T_809 = _T_805 & _T_808;
  assign _T_810 = _T_809[6:4];
  assign _T_811 = _T_809[3:0];
  assign _T_813 = _T_810 != 3'h0;
  assign _GEN_51 = {{1'd0}, _T_810};
  assign _T_814 = _GEN_51 | _T_811;
  assign _T_815 = _T_814[3:2];
  assign _T_816 = _T_814[1:0];
  assign _T_818 = _T_815 != 2'h0;
  assign _T_819 = _T_815 | _T_816;
  assign _T_820 = _T_819[1];
  assign _T_821 = {_T_818,_T_820};
  assign _T_822 = {_T_813,_T_821};
  assign _T_823 = io_out_2_d_ready & io_out_2_d_valid;
  assign _GEN_52 = {{3'd0}, _T_800};
  assign _T_824 = _T_763 - _GEN_52;
  assign _T_825 = $unsigned(_T_824);
  assign _T_826 = _T_825[3:0];
  assign _T_827 = _T_771 ? _T_769 : _T_826;
  assign _T_828 = io_out_2_d_bits_source[4];
  assign _GEN_16 = _T_771 ? _T_822 : _T_765;
  assign _GEN_17 = _T_771 ? _T_828 : _T_768;
  assign _GEN_18 = _T_823 ? _T_827 : _T_763;
  assign _GEN_19 = _T_823 ? _GEN_16 : _T_765;
  assign _GEN_20 = _T_823 ? _GEN_17 : _T_768;
  assign _T_830 = _T_783 == 1'h0;
  assign _T_832 = _T_773 == 1'h0;
  assign _T_833 = _T_830 & _T_832;
  assign _T_834 = io_in_2_d_ready | _T_833;
  assign _T_836 = _T_833 == 1'h0;
  assign _T_837 = io_out_2_d_valid & _T_836;
  assign _T_838 = io_out_2_d_bits_source[9:5];
  assign _T_843 = _T_842 | io_out_2_d_bits_error;
  assign _T_846 = _T_833 ? _T_843 : 1'h0;
  assign _GEN_21 = _T_823 ? _T_846 : _T_842;
  assign Repeater_2_clock = clock;
  assign Repeater_2_reset = reset;
  assign Repeater_2_io_repeat = _T_932;
  assign Repeater_2_io_enq_valid = io_in_2_a_valid;
  assign Repeater_2_io_enq_bits_opcode = io_in_2_a_bits_opcode;
  assign Repeater_2_io_enq_bits_size = io_in_2_a_bits_size;
  assign Repeater_2_io_enq_bits_source = io_in_2_a_bits_source;
  assign Repeater_2_io_enq_bits_address = io_in_2_a_bits_address;
  assign Repeater_2_io_enq_bits_mask = io_in_2_a_bits_mask;
  assign Repeater_2_io_deq_ready = io_out_2_a_ready;
  assign _T_883 = Repeater_2_io_deq_bits_size > 3'h2;
  assign _T_884 = _T_883 ? 3'h2 : Repeater_2_io_deq_bits_size;
  assign _T_887 = 13'h3f << Repeater_2_io_deq_bits_size;
  assign _T_888 = _T_887[5:0];
  assign _T_889 = ~ _T_888;
  assign _T_892 = 9'h3 << _T_884;
  assign _T_893 = _T_892[1:0];
  assign _T_894 = ~ _T_893;
  assign _T_895 = Repeater_2_io_deq_bits_opcode[2];
  assign _T_897 = _T_895 == 1'h0;
  assign _T_904 = _T_902 == 4'h0;
  assign _T_905 = _T_889[5:2];
  assign _T_907 = _T_902 - 4'h1;
  assign _T_908 = $unsigned(_T_907);
  assign _T_909 = _T_908[3:0];
  assign _T_910 = _T_904 ? _T_905 : _T_909;
  assign _T_911 = ~ _T_910;
  assign _T_914 = ~ _T_911;
  assign _GEN_22 = _T_904 ? _T_768 : _T_923;
  assign _T_926 = _GEN_22 == 1'h0;
  assign _T_927 = io_out_2_a_ready & io_out_2_a_valid;
  assign _GEN_23 = _T_927 ? _T_914 : _T_902;
  assign _T_929 = _T_897 == 1'h0;
  assign _T_931 = _T_914 != 4'h0;
  assign _T_932 = _T_929 & _T_931;
  assign _GEN_53 = {{2'd0}, _T_910};
  assign _T_933 = _GEN_53 << 2;
  assign _T_934 = ~ _T_889;
  assign _T_935 = _T_933 | _T_934;
  assign _GEN_54 = {{4'd0}, _T_894};
  assign _T_936 = _T_935 | _GEN_54;
  assign _T_938 = _T_936 | 6'h3;
  assign _T_939 = ~ _T_938;
  assign _GEN_55 = {{6'd0}, _T_939};
  assign _T_940 = Repeater_2_io_deq_bits_address | _GEN_55;
  assign _T_941 = {Repeater_2_io_deq_bits_source,_T_926};
  assign _T_942 = {_T_941,_T_914};
  assign _T_944 = Repeater_2_io_full == 1'h0;
  assign _T_947 = _T_944 | _T_929;
  assign _T_948 = _T_947 | reset;
  assign _T_950 = _T_948 == 1'h0;
  assign _T_954 = Repeater_2_io_deq_bits_mask == 4'hf;
  assign _T_955 = _T_944 | _T_954;
  assign _T_956 = _T_955 | reset;
  assign _T_958 = _T_956 == 1'h0;
  assign _T_959 = Repeater_2_io_full ? 4'hf : io_in_2_a_bits_mask;
  assign _T_974 = io_out_3_d_bits_source[3:0];
  assign _T_976 = _T_968 == 4'h0;
  assign _T_985 = 5'h3 << io_out_3_d_bits_size;
  assign _T_986 = _T_985[1:0];
  assign _T_987 = ~ _T_986;
  assign _GEN_56 = {{2'd0}, _T_974};
  assign _T_1007 = _GEN_56 << 2;
  assign _GEN_57 = {{4'd0}, _T_987};
  assign _T_1008 = _T_1007 | _GEN_57;
  assign _GEN_58 = {{1'd0}, _T_1008};
  assign _T_1009 = _GEN_58 << 1;
  assign _T_1011 = _T_1009 | 7'h1;
  assign _T_1013 = {1'h0,_T_1008};
  assign _T_1014 = ~ _T_1013;
  assign _T_1015 = _T_1011 & _T_1014;
  assign _T_1016 = _T_1015[6:4];
  assign _T_1017 = _T_1015[3:0];
  assign _T_1019 = _T_1016 != 3'h0;
  assign _GEN_59 = {{1'd0}, _T_1016};
  assign _T_1020 = _GEN_59 | _T_1017;
  assign _T_1021 = _T_1020[3:2];
  assign _T_1022 = _T_1020[1:0];
  assign _T_1024 = _T_1021 != 2'h0;
  assign _T_1025 = _T_1021 | _T_1022;
  assign _T_1026 = _T_1025[1];
  assign _T_1027 = {_T_1024,_T_1026};
  assign _T_1028 = {_T_1019,_T_1027};
  assign _T_1029 = io_out_3_d_ready & io_out_3_d_valid;
  assign _T_1030 = _T_968 - 4'h1;
  assign _T_1031 = $unsigned(_T_1030);
  assign _T_1032 = _T_1031[3:0];
  assign _T_1033 = _T_976 ? _T_974 : _T_1032;
  assign _T_1034 = io_out_3_d_bits_source[4];
  assign _GEN_24 = _T_976 ? _T_1028 : _T_970;
  assign _GEN_25 = _T_976 ? _T_1034 : _T_973;
  assign _GEN_26 = _T_1029 ? _T_1033 : _T_968;
  assign _GEN_27 = _T_1029 ? _GEN_24 : _T_970;
  assign _GEN_28 = _T_1029 ? _GEN_25 : _T_973;
  assign _T_1044 = io_out_3_d_bits_source[9:5];
  assign _T_1049 = _T_1048 | io_out_3_d_bits_error;
  assign _GEN_29 = _T_1029 ? 1'h0 : _T_1048;
  assign Repeater_3_clock = clock;
  assign Repeater_3_reset = reset;
  assign Repeater_3_io_repeat = _T_1136;
  assign Repeater_3_io_enq_valid = io_in_3_a_valid;
  assign Repeater_3_io_enq_bits_opcode = io_in_3_a_bits_opcode;
  assign Repeater_3_io_enq_bits_size = io_in_3_a_bits_size;
  assign Repeater_3_io_enq_bits_source = io_in_3_a_bits_source;
  assign Repeater_3_io_enq_bits_address = io_in_3_a_bits_address;
  assign Repeater_3_io_enq_bits_mask = io_in_3_a_bits_mask;
  assign Repeater_3_io_deq_ready = io_out_3_a_ready;
  assign _T_1087 = Repeater_3_io_deq_bits_size > 3'h2;
  assign _T_1088 = _T_1087 ? 3'h2 : Repeater_3_io_deq_bits_size;
  assign _T_1091 = 13'h3f << Repeater_3_io_deq_bits_size;
  assign _T_1092 = _T_1091[5:0];
  assign _T_1093 = ~ _T_1092;
  assign _T_1096 = 9'h3 << _T_1088;
  assign _T_1097 = _T_1096[1:0];
  assign _T_1098 = ~ _T_1097;
  assign _T_1099 = Repeater_3_io_deq_bits_opcode[2];
  assign _T_1101 = _T_1099 == 1'h0;
  assign _T_1108 = _T_1106 == 4'h0;
  assign _T_1109 = _T_1093[5:2];
  assign _T_1111 = _T_1106 - 4'h1;
  assign _T_1112 = $unsigned(_T_1111);
  assign _T_1113 = _T_1112[3:0];
  assign _T_1114 = _T_1108 ? _T_1109 : _T_1113;
  assign _T_1115 = ~ _T_1114;
  assign _T_1118 = ~ _T_1115;
  assign _GEN_30 = _T_1108 ? _T_973 : _T_1127;
  assign _T_1130 = _GEN_30 == 1'h0;
  assign _T_1131 = io_out_3_a_ready & io_out_3_a_valid;
  assign _GEN_31 = _T_1131 ? _T_1118 : _T_1106;
  assign _T_1133 = _T_1101 == 1'h0;
  assign _T_1135 = _T_1118 != 4'h0;
  assign _T_1136 = _T_1133 & _T_1135;
  assign _GEN_60 = {{2'd0}, _T_1114};
  assign _T_1137 = _GEN_60 << 2;
  assign _T_1138 = ~ _T_1093;
  assign _T_1139 = _T_1137 | _T_1138;
  assign _GEN_61 = {{4'd0}, _T_1098};
  assign _T_1140 = _T_1139 | _GEN_61;
  assign _T_1142 = _T_1140 | 6'h3;
  assign _T_1143 = ~ _T_1142;
  assign _GEN_62 = {{11'd0}, _T_1143};
  assign _T_1144 = Repeater_3_io_deq_bits_address | _GEN_62;
  assign _T_1145 = {Repeater_3_io_deq_bits_source,_T_1130};
  assign _T_1146 = {_T_1145,_T_1118};
  assign _T_1148 = Repeater_3_io_full == 1'h0;
  assign _T_1151 = _T_1148 | _T_1133;
  assign _T_1152 = _T_1151 | reset;
  assign _T_1154 = _T_1152 == 1'h0;
  assign _T_1158 = Repeater_3_io_deq_bits_mask == 4'hf;
  assign _T_1159 = _T_1148 | _T_1158;
  assign _T_1160 = _T_1159 | reset;
  assign _T_1162 = _T_1160 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_353 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_355 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_358 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_432 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_492 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_513 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_558 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_560 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_563 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_637 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_697 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_718 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_763 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_765 = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_768 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_842 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_902 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_923 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_968 = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_970 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_973 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_1048 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_1106 = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_1127 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_353 <= 4'h0;
    end else begin
      if (_T_413) begin
        if (_T_361) begin
          _T_353 <= _T_359;
        end else begin
          _T_353 <= _T_416;
        end
      end
    end
    if (_T_413) begin
      if (_T_361) begin
        _T_355 <= _T_412;
      end
    end
    if (reset) begin
      _T_358 <= 1'h0;
    end else begin
      if (_T_413) begin
        if (_T_361) begin
          _T_358 <= _T_418;
        end
      end
    end
    if (reset) begin
      _T_432 <= 1'h0;
    end else begin
      if (_T_413) begin
        if (_T_423) begin
          _T_432 <= _T_433;
        end else begin
          _T_432 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_492 <= 4'h0;
    end else begin
      if (_T_517) begin
        _T_492 <= _T_504;
      end
    end
    if (_T_494) begin
      _T_513 <= _T_358;
    end
    if (reset) begin
      _T_558 <= 4'h0;
    end else begin
      if (_T_618) begin
        if (_T_566) begin
          _T_558 <= _T_564;
        end else begin
          _T_558 <= _T_621;
        end
      end
    end
    if (_T_618) begin
      if (_T_566) begin
        _T_560 <= _T_617;
      end
    end
    if (reset) begin
      _T_563 <= 1'h0;
    end else begin
      if (_T_618) begin
        if (_T_566) begin
          _T_563 <= _T_623;
        end
      end
    end
    if (reset) begin
      _T_637 <= 1'h0;
    end else begin
      if (_T_618) begin
        if (_T_628) begin
          _T_637 <= _T_638;
        end else begin
          _T_637 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_697 <= 4'h0;
    end else begin
      if (_T_722) begin
        _T_697 <= _T_709;
      end
    end
    if (_T_699) begin
      _T_718 <= _T_563;
    end
    if (reset) begin
      _T_763 <= 4'h0;
    end else begin
      if (_T_823) begin
        if (_T_771) begin
          _T_763 <= _T_769;
        end else begin
          _T_763 <= _T_826;
        end
      end
    end
    if (_T_823) begin
      if (_T_771) begin
        _T_765 <= _T_822;
      end
    end
    if (reset) begin
      _T_768 <= 1'h0;
    end else begin
      if (_T_823) begin
        if (_T_771) begin
          _T_768 <= _T_828;
        end
      end
    end
    if (reset) begin
      _T_842 <= 1'h0;
    end else begin
      if (_T_823) begin
        if (_T_833) begin
          _T_842 <= _T_843;
        end else begin
          _T_842 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_902 <= 4'h0;
    end else begin
      if (_T_927) begin
        _T_902 <= _T_914;
      end
    end
    if (_T_904) begin
      _T_923 <= _T_768;
    end
    if (reset) begin
      _T_968 <= 4'h0;
    end else begin
      if (_T_1029) begin
        if (_T_976) begin
          _T_968 <= _T_974;
        end else begin
          _T_968 <= _T_1032;
        end
      end
    end
    if (_T_1029) begin
      if (_T_976) begin
        _T_970 <= _T_1028;
      end
    end
    if (reset) begin
      _T_973 <= 1'h0;
    end else begin
      if (_T_1029) begin
        if (_T_976) begin
          _T_973 <= _T_1034;
        end
      end
    end
    if (reset) begin
      _T_1048 <= 1'h0;
    end else begin
      if (_T_1029) begin
        _T_1048 <= 1'h0;
      end
    end
    if (reset) begin
      _T_1106 <= 4'h0;
    end else begin
      if (_T_1131) begin
        _T_1106 <= _T_1118;
      end
    end
    if (_T_1108) begin
      _T_1127 <= _T_973;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:174 assert (!out.d.valid || (acknum_fragment & acknum_size) === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_540) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:273 assert (!repeater.io.full || !aHasData)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_540) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_548) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:276 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_548) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:174 assert (!out.d.valid || (acknum_fragment & acknum_size) === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_745) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:273 assert (!repeater.io.full || !aHasData)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_745) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_753) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:276 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_753) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:174 assert (!out.d.valid || (acknum_fragment & acknum_size) === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_950) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:273 assert (!repeater.io.full || !aHasData)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_950) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_958) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:276 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_958) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:174 assert (!out.d.valid || (acknum_fragment & acknum_size) === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1154) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:273 assert (!repeater.io.full || !aHasData)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1154) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1162) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:276 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1162) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module TLAtomicAutomata(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [2:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [2:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  reg [1:0] _T_108_0_state;
  reg [31:0] _RAND_0;
  reg [2:0] _T_119_0_bits_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] _T_119_0_bits_param;
  reg [31:0] _RAND_2;
  reg [2:0] _T_119_0_bits_size;
  reg [31:0] _RAND_3;
  reg [4:0] _T_119_0_bits_source;
  reg [31:0] _RAND_4;
  reg [31:0] _T_119_0_bits_address;
  reg [31:0] _RAND_5;
  reg [3:0] _T_119_0_bits_mask;
  reg [31:0] _RAND_6;
  reg [31:0] _T_119_0_bits_data;
  reg [31:0] _RAND_7;
  reg [1:0] _T_119_0_fifoId;
  reg [31:0] _RAND_8;
  reg [3:0] _T_119_0_lut;
  reg [31:0] _RAND_9;
  reg [31:0] _T_126_0_data;
  reg [31:0] _RAND_10;
  wire  _T_130;
  wire  _T_131;
  wire  _T_132;
  wire  _T_134;
  wire  _T_135;
  wire  _T_139;
  wire [31:0] _T_142;
  wire [32:0] _T_143;
  wire [32:0] _T_145;
  wire [32:0] _T_146;
  wire  _T_148;
  wire  _T_149;
  wire [32:0] _T_155;
  wire  _T_197;
  wire  _T_199;
  wire  _T_201;
  wire  _T_202;
  wire [32:0] _T_212;
  wire [32:0] _T_213;
  wire  _T_215;
  wire [31:0] _T_218;
  wire [32:0] _T_219;
  wire [32:0] _T_221;
  wire [32:0] _T_222;
  wire  _T_224;
  wire [32:0] _T_230;
  wire [32:0] _T_231;
  wire  _T_233;
  wire [1:0] _T_255;
  wire [1:0] _T_259;
  wire [1:0] _GEN_31;
  wire [1:0] _T_262;
  wire [1:0] _T_263;
  wire  _T_267;
  wire  _T_268;
  wire  _T_274;
  wire  _T_275;
  wire [1:0] _T_276;
  wire  _T_277;
  wire  _T_278;
  wire [1:0] _T_279;
  wire  _T_280;
  wire  _T_281;
  wire [1:0] _T_282;
  wire  _T_283;
  wire  _T_284;
  wire [1:0] _T_285;
  wire  _T_286;
  wire  _T_287;
  wire [1:0] _T_288;
  wire  _T_289;
  wire  _T_290;
  wire [1:0] _T_291;
  wire  _T_292;
  wire  _T_293;
  wire [1:0] _T_294;
  wire  _T_295;
  wire  _T_296;
  wire [1:0] _T_297;
  wire  _T_298;
  wire  _T_299;
  wire [1:0] _T_300;
  wire  _T_301;
  wire  _T_302;
  wire [1:0] _T_303;
  wire  _T_304;
  wire  _T_305;
  wire [1:0] _T_306;
  wire  _T_307;
  wire  _T_308;
  wire [1:0] _T_309;
  wire  _T_310;
  wire  _T_311;
  wire [1:0] _T_312;
  wire  _T_313;
  wire  _T_314;
  wire [1:0] _T_315;
  wire  _T_316;
  wire  _T_317;
  wire [1:0] _T_318;
  wire  _T_319;
  wire  _T_320;
  wire [1:0] _T_321;
  wire  _T_322;
  wire  _T_323;
  wire [1:0] _T_324;
  wire  _T_325;
  wire  _T_326;
  wire [1:0] _T_327;
  wire  _T_328;
  wire  _T_329;
  wire [1:0] _T_330;
  wire  _T_331;
  wire  _T_332;
  wire [1:0] _T_333;
  wire  _T_334;
  wire  _T_335;
  wire [1:0] _T_336;
  wire  _T_337;
  wire  _T_338;
  wire [1:0] _T_339;
  wire  _T_340;
  wire  _T_341;
  wire [1:0] _T_342;
  wire  _T_343;
  wire  _T_344;
  wire [1:0] _T_345;
  wire  _T_346;
  wire  _T_347;
  wire [1:0] _T_348;
  wire  _T_349;
  wire  _T_350;
  wire [1:0] _T_351;
  wire  _T_352;
  wire  _T_353;
  wire [1:0] _T_354;
  wire  _T_355;
  wire  _T_356;
  wire [1:0] _T_357;
  wire  _T_358;
  wire  _T_359;
  wire [1:0] _T_360;
  wire  _T_361;
  wire  _T_362;
  wire [1:0] _T_363;
  wire  _T_364;
  wire  _T_365;
  wire [1:0] _T_366;
  wire  _T_367;
  wire  _T_368;
  wire [1:0] _T_369;
  wire [3:0] _T_370;
  wire  _T_371;
  wire [3:0] _T_372;
  wire  _T_373;
  wire [3:0] _T_374;
  wire  _T_375;
  wire [3:0] _T_376;
  wire  _T_377;
  wire [3:0] _T_378;
  wire  _T_379;
  wire [3:0] _T_380;
  wire  _T_381;
  wire [3:0] _T_382;
  wire  _T_383;
  wire [3:0] _T_384;
  wire  _T_385;
  wire [3:0] _T_386;
  wire  _T_387;
  wire [3:0] _T_388;
  wire  _T_389;
  wire [3:0] _T_390;
  wire  _T_391;
  wire [3:0] _T_392;
  wire  _T_393;
  wire [3:0] _T_394;
  wire  _T_395;
  wire [3:0] _T_396;
  wire  _T_397;
  wire [3:0] _T_398;
  wire  _T_399;
  wire [3:0] _T_400;
  wire  _T_401;
  wire [3:0] _T_402;
  wire  _T_403;
  wire [3:0] _T_404;
  wire  _T_405;
  wire [3:0] _T_406;
  wire  _T_407;
  wire [3:0] _T_408;
  wire  _T_409;
  wire [3:0] _T_410;
  wire  _T_411;
  wire [3:0] _T_412;
  wire  _T_413;
  wire [3:0] _T_414;
  wire  _T_415;
  wire [3:0] _T_416;
  wire  _T_417;
  wire [3:0] _T_418;
  wire  _T_419;
  wire [3:0] _T_420;
  wire  _T_421;
  wire [3:0] _T_422;
  wire  _T_423;
  wire [3:0] _T_424;
  wire  _T_425;
  wire [3:0] _T_426;
  wire  _T_427;
  wire [3:0] _T_428;
  wire  _T_429;
  wire [3:0] _T_430;
  wire  _T_431;
  wire [3:0] _T_432;
  wire  _T_433;
  wire [1:0] _T_434;
  wire [1:0] _T_435;
  wire [3:0] _T_436;
  wire [1:0] _T_437;
  wire [1:0] _T_438;
  wire [3:0] _T_439;
  wire [7:0] _T_440;
  wire [1:0] _T_441;
  wire [1:0] _T_442;
  wire [3:0] _T_443;
  wire [1:0] _T_444;
  wire [1:0] _T_445;
  wire [3:0] _T_446;
  wire [7:0] _T_447;
  wire [15:0] _T_448;
  wire [1:0] _T_449;
  wire [1:0] _T_450;
  wire [3:0] _T_451;
  wire [1:0] _T_452;
  wire [1:0] _T_453;
  wire [3:0] _T_454;
  wire [7:0] _T_455;
  wire [1:0] _T_456;
  wire [1:0] _T_457;
  wire [3:0] _T_458;
  wire [1:0] _T_459;
  wire [1:0] _T_460;
  wire [3:0] _T_461;
  wire [7:0] _T_462;
  wire [15:0] _T_463;
  wire [31:0] _T_464;
  wire  _T_465;
  wire  _T_466;
  wire  _T_467;
  wire [3:0] _T_468;
  wire [2:0] _T_469;
  wire [3:0] _GEN_32;
  wire [3:0] _T_470;
  wire [3:0] _T_471;
  wire [1:0] _T_476;
  wire [1:0] _T_477;
  wire [3:0] _T_478;
  wire [1:0] _T_483;
  wire [1:0] _T_484;
  wire [3:0] _T_485;
  wire [3:0] _T_486;
  wire [4:0] _GEN_33;
  wire [4:0] _T_487;
  wire [3:0] _T_488;
  wire [3:0] _T_489;
  wire [4:0] _GEN_34;
  wire [4:0] _T_490;
  wire [3:0] _T_491;
  wire [4:0] _GEN_35;
  wire [4:0] _T_492;
  wire [3:0] _T_493;
  wire [3:0] _T_494;
  wire [5:0] _GEN_36;
  wire [5:0] _T_495;
  wire [3:0] _T_496;
  wire [3:0] _T_497;
  wire  _T_499;
  wire  _T_500;
  wire  _T_501;
  wire  _T_502;
  wire [7:0] _T_506;
  wire [7:0] _T_510;
  wire [7:0] _T_514;
  wire [7:0] _T_518;
  wire [15:0] _T_519;
  wire [15:0] _T_520;
  wire [31:0] _T_521;
  wire [4:0] _GEN_37;
  wire [4:0] _T_522;
  wire [3:0] _T_523;
  wire [3:0] _T_524;
  wire [5:0] _GEN_38;
  wire [5:0] _T_525;
  wire [3:0] _T_526;
  wire [3:0] _T_527;
  wire  _T_529;
  wire  _T_530;
  wire  _T_531;
  wire  _T_532;
  wire [7:0] _T_536;
  wire [7:0] _T_540;
  wire [7:0] _T_544;
  wire [7:0] _T_548;
  wire [15:0] _T_549;
  wire [15:0] _T_550;
  wire [31:0] _T_551;
  wire  _T_552;
  wire  _T_553;
  wire  _T_554;
  wire  _T_555;
  wire [7:0] _T_559;
  wire [7:0] _T_563;
  wire [7:0] _T_567;
  wire [7:0] _T_571;
  wire [15:0] _T_572;
  wire [15:0] _T_573;
  wire [31:0] _T_574;
  wire [31:0] _T_575;
  wire [31:0] _T_576;
  wire [31:0] _T_577;
  wire [31:0] _T_578;
  wire [31:0] _T_579;
  wire [31:0] _T_580;
  wire [32:0] _T_581;
  wire [31:0] _T_582;
  wire  _T_583;
  wire  _T_584;
  wire  _T_586;
  wire  _T_587;
  wire  _T_588;
  wire  _T_590;
  wire  _T_591;
  wire  _T_592;
  wire [31:0] _T_593;
  wire [31:0] _T_594;
  wire  _T_595;
  wire [31:0] _T_596;
  wire  _T_602;
  wire  _T_603;
  wire  _T_604;
  wire  _T_605;
  wire  _T_606;
  wire  _T_608;
  wire [2:0] _GEN_0;
  wire [2:0] _GEN_1;
  wire  _T_659;
  wire [1:0] _T_661;
  wire [1:0] _T_664;
  wire  _T_666;
  wire  _T_668;
  wire  _T_669;
  wire  _T_671;
  wire  _T_673;
  wire  _T_674;
  wire  _T_676;
  wire  _T_677;
  wire  _T_678;
  wire  _T_679;
  wire  _T_681;
  wire  _T_682;
  wire  _T_683;
  wire  _T_684;
  wire  _T_685;
  wire  _T_686;
  wire  _T_687;
  wire  _T_688;
  wire  _T_689;
  wire  _T_690;
  wire  _T_691;
  wire  _T_692;
  wire  _T_693;
  wire [1:0] _T_694;
  wire [1:0] _T_695;
  wire [3:0] _T_696;
  wire [12:0] _T_700;
  wire [5:0] _T_701;
  wire [5:0] _T_702;
  wire [3:0] _T_703;
  wire  _T_704;
  wire  _T_706;
  wire [3:0] _T_708;
  reg [3:0] _T_711;
  reg [31:0] _RAND_11;
  wire  _T_713;
  wire  _T_714;
  wire [1:0] _T_715;
  wire [2:0] _GEN_39;
  wire [2:0] _T_716;
  wire [1:0] _T_717;
  wire [1:0] _T_718;
  wire [2:0] _GEN_40;
  wire [2:0] _T_720;
  wire [1:0] _T_721;
  wire [1:0] _T_722;
  wire  _T_723;
  wire  _T_724;
  wire  _T_732;
  wire  _T_733;
  wire  _T_743;
  wire  _T_747;
  wire  _T_752;
  wire  _T_753;
  wire  _T_755;
  wire  _T_757;
  wire  _T_758;
  wire  _T_760;
  wire  _T_762;
  wire  _T_763;
  wire  _T_765;
  wire [3:0] _T_769;
  wire  _T_771;
  wire [3:0] _GEN_41;
  wire [4:0] _T_772;
  wire [4:0] _T_773;
  wire [3:0] _T_774;
  wire [3:0] _T_775;
  reg  _T_793_0;
  reg [31:0] _RAND_12;
  reg  _T_793_1;
  reg [31:0] _RAND_13;
  wire  _T_804_0;
  wire  _T_804_1;
  wire  _T_812_0;
  wire  _T_812_1;
  wire  _T_820;
  wire  _T_821;
  wire  _T_825;
  wire  _T_827;
  wire  _T_828;
  wire  _T_831;
  wire [35:0] _T_833;
  wire [67:0] _T_834;
  wire [7:0] _T_835;
  wire [13:0] _T_837;
  wire [81:0] _T_838;
  wire [81:0] _T_840;
  wire [35:0] _T_841;
  wire [67:0] _T_842;
  wire [7:0] _T_843;
  wire [5:0] _T_844;
  wire [13:0] _T_845;
  wire [81:0] _T_846;
  wire [81:0] _T_848;
  wire [81:0] _T_849;
  wire [31:0] _T_854;
  wire [3:0] _T_855;
  wire [31:0] _T_856;
  wire [4:0] _T_857;
  wire [2:0] _T_858;
  wire [2:0] _T_859;
  wire [2:0] _T_860;
  wire  _T_861;
  wire  _T_864;
  wire [1:0] _T_865;
  wire [2:0] _GEN_42;
  wire  _T_875;
  wire [3:0] _T_876;
  wire  _T_877;
  wire [3:0] _T_878;
  wire  _T_879;
  wire [3:0] _T_880;
  wire  _T_881;
  wire [3:0] _T_882;
  wire [1:0] _GEN_2;
  wire [2:0] _GEN_3;
  wire [2:0] _GEN_4;
  wire [2:0] _GEN_5;
  wire [4:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [3:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [3:0] _GEN_10;
  wire [1:0] _GEN_11;
  wire [1:0] _GEN_12;
  wire [2:0] _GEN_13;
  wire [2:0] _GEN_14;
  wire [2:0] _GEN_15;
  wire [4:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [3:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [3:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire  _T_883;
  wire [1:0] _GEN_22;
  wire [1:0] _GEN_23;
  wire  _T_884;
  wire [12:0] _T_887;
  wire [5:0] _T_888;
  wire [5:0] _T_889;
  wire [3:0] _T_890;
  wire  _T_891;
  wire [3:0] _T_893;
  reg [3:0] _T_896;
  reg [31:0] _RAND_14;
  wire [4:0] _T_898;
  wire [4:0] _T_899;
  wire [3:0] _T_900;
  wire  _T_902;
  wire [3:0] _T_911;
  wire [3:0] _GEN_24;
  wire  _T_912;
  wire  _T_913;
  wire  _T_918;
  wire  _T_920;
  wire  _T_922;
  wire  _T_923;
  wire [31:0] _GEN_25;
  wire [1:0] _T_924;
  wire [1:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire [1:0] _GEN_28;
  wire  _T_925;
  wire  _T_926;
  wire  _T_927;
  wire  _T_928;
  wire  _T_930;
  wire  _T_931;
  wire  _T_932;
  wire [2:0] _GEN_29;
  wire [31:0] _GEN_30;
  assign io_in_0_a_ready = _T_605;
  assign io_in_0_d_valid = _T_931;
  assign io_in_0_d_bits_opcode = _GEN_29;
  assign io_in_0_d_bits_param = io_out_0_d_bits_param;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_in_0_d_bits_sink = io_out_0_d_bits_sink;
  assign io_in_0_d_bits_data = _GEN_30;
  assign io_in_0_d_bits_error = io_out_0_d_bits_error;
  assign io_out_0_a_valid = _T_831;
  assign io_out_0_a_bits_opcode = _T_860;
  assign io_out_0_a_bits_param = _T_859;
  assign io_out_0_a_bits_size = _T_858;
  assign io_out_0_a_bits_source = _T_857;
  assign io_out_0_a_bits_address = _T_856;
  assign io_out_0_a_bits_mask = _T_855;
  assign io_out_0_a_bits_data = _T_854;
  assign io_out_0_d_ready = _T_932;
  assign _T_130 = _T_108_0_state == 2'h0;
  assign _T_131 = _T_108_0_state == 2'h2;
  assign _T_132 = _T_108_0_state == 2'h3;
  assign _T_134 = _T_132 | _T_131;
  assign _T_135 = _T_108_0_state != 2'h0;
  assign _T_139 = 3'h2 == io_in_0_a_bits_size;
  assign _T_142 = io_in_0_a_bits_address ^ 32'h80000000;
  assign _T_143 = {1'b0,$signed(_T_142)};
  assign _T_145 = $signed(_T_143) & $signed(33'sh80000000);
  assign _T_146 = $signed(_T_145);
  assign _T_148 = $signed(_T_146) == $signed(33'sh0);
  assign _T_149 = _T_139 & _T_148;
  assign _T_155 = {1'b0,$signed(io_in_0_a_bits_address)};
  assign _T_197 = io_in_0_a_bits_opcode == 3'h3;
  assign _T_199 = io_in_0_a_bits_opcode == 3'h2;
  assign _T_201 = _T_199 ? _T_149 : 1'h1;
  assign _T_202 = _T_197 ? _T_149 : _T_201;
  assign _T_212 = $signed(_T_155) & $signed(33'sh86010000);
  assign _T_213 = $signed(_T_212);
  assign _T_215 = $signed(_T_213) == $signed(33'sh0);
  assign _T_218 = io_in_0_a_bits_address ^ 32'h2000000;
  assign _T_219 = {1'b0,$signed(_T_218)};
  assign _T_221 = $signed(_T_219) & $signed(33'sh86010000);
  assign _T_222 = $signed(_T_221);
  assign _T_224 = $signed(_T_222) == $signed(33'sh0);
  assign _T_230 = $signed(_T_143) & $signed(33'sh86010000);
  assign _T_231 = $signed(_T_230);
  assign _T_233 = $signed(_T_231) == $signed(33'sh0);
  assign _T_255 = _T_215 ? 2'h2 : 2'h0;
  assign _T_259 = _T_233 ? 2'h3 : 2'h0;
  assign _GEN_31 = {{1'd0}, _T_224};
  assign _T_262 = _T_255 | _GEN_31;
  assign _T_263 = _T_262 | _T_259;
  assign _T_267 = _T_119_0_fifoId == _T_263;
  assign _T_268 = _T_134 & _T_267;
  assign _T_274 = _T_119_0_bits_data[0];
  assign _T_275 = _T_126_0_data[0];
  assign _T_276 = {_T_274,_T_275};
  assign _T_277 = _T_119_0_bits_data[1];
  assign _T_278 = _T_126_0_data[1];
  assign _T_279 = {_T_277,_T_278};
  assign _T_280 = _T_119_0_bits_data[2];
  assign _T_281 = _T_126_0_data[2];
  assign _T_282 = {_T_280,_T_281};
  assign _T_283 = _T_119_0_bits_data[3];
  assign _T_284 = _T_126_0_data[3];
  assign _T_285 = {_T_283,_T_284};
  assign _T_286 = _T_119_0_bits_data[4];
  assign _T_287 = _T_126_0_data[4];
  assign _T_288 = {_T_286,_T_287};
  assign _T_289 = _T_119_0_bits_data[5];
  assign _T_290 = _T_126_0_data[5];
  assign _T_291 = {_T_289,_T_290};
  assign _T_292 = _T_119_0_bits_data[6];
  assign _T_293 = _T_126_0_data[6];
  assign _T_294 = {_T_292,_T_293};
  assign _T_295 = _T_119_0_bits_data[7];
  assign _T_296 = _T_126_0_data[7];
  assign _T_297 = {_T_295,_T_296};
  assign _T_298 = _T_119_0_bits_data[8];
  assign _T_299 = _T_126_0_data[8];
  assign _T_300 = {_T_298,_T_299};
  assign _T_301 = _T_119_0_bits_data[9];
  assign _T_302 = _T_126_0_data[9];
  assign _T_303 = {_T_301,_T_302};
  assign _T_304 = _T_119_0_bits_data[10];
  assign _T_305 = _T_126_0_data[10];
  assign _T_306 = {_T_304,_T_305};
  assign _T_307 = _T_119_0_bits_data[11];
  assign _T_308 = _T_126_0_data[11];
  assign _T_309 = {_T_307,_T_308};
  assign _T_310 = _T_119_0_bits_data[12];
  assign _T_311 = _T_126_0_data[12];
  assign _T_312 = {_T_310,_T_311};
  assign _T_313 = _T_119_0_bits_data[13];
  assign _T_314 = _T_126_0_data[13];
  assign _T_315 = {_T_313,_T_314};
  assign _T_316 = _T_119_0_bits_data[14];
  assign _T_317 = _T_126_0_data[14];
  assign _T_318 = {_T_316,_T_317};
  assign _T_319 = _T_119_0_bits_data[15];
  assign _T_320 = _T_126_0_data[15];
  assign _T_321 = {_T_319,_T_320};
  assign _T_322 = _T_119_0_bits_data[16];
  assign _T_323 = _T_126_0_data[16];
  assign _T_324 = {_T_322,_T_323};
  assign _T_325 = _T_119_0_bits_data[17];
  assign _T_326 = _T_126_0_data[17];
  assign _T_327 = {_T_325,_T_326};
  assign _T_328 = _T_119_0_bits_data[18];
  assign _T_329 = _T_126_0_data[18];
  assign _T_330 = {_T_328,_T_329};
  assign _T_331 = _T_119_0_bits_data[19];
  assign _T_332 = _T_126_0_data[19];
  assign _T_333 = {_T_331,_T_332};
  assign _T_334 = _T_119_0_bits_data[20];
  assign _T_335 = _T_126_0_data[20];
  assign _T_336 = {_T_334,_T_335};
  assign _T_337 = _T_119_0_bits_data[21];
  assign _T_338 = _T_126_0_data[21];
  assign _T_339 = {_T_337,_T_338};
  assign _T_340 = _T_119_0_bits_data[22];
  assign _T_341 = _T_126_0_data[22];
  assign _T_342 = {_T_340,_T_341};
  assign _T_343 = _T_119_0_bits_data[23];
  assign _T_344 = _T_126_0_data[23];
  assign _T_345 = {_T_343,_T_344};
  assign _T_346 = _T_119_0_bits_data[24];
  assign _T_347 = _T_126_0_data[24];
  assign _T_348 = {_T_346,_T_347};
  assign _T_349 = _T_119_0_bits_data[25];
  assign _T_350 = _T_126_0_data[25];
  assign _T_351 = {_T_349,_T_350};
  assign _T_352 = _T_119_0_bits_data[26];
  assign _T_353 = _T_126_0_data[26];
  assign _T_354 = {_T_352,_T_353};
  assign _T_355 = _T_119_0_bits_data[27];
  assign _T_356 = _T_126_0_data[27];
  assign _T_357 = {_T_355,_T_356};
  assign _T_358 = _T_119_0_bits_data[28];
  assign _T_359 = _T_126_0_data[28];
  assign _T_360 = {_T_358,_T_359};
  assign _T_361 = _T_119_0_bits_data[29];
  assign _T_362 = _T_126_0_data[29];
  assign _T_363 = {_T_361,_T_362};
  assign _T_364 = _T_119_0_bits_data[30];
  assign _T_365 = _T_126_0_data[30];
  assign _T_366 = {_T_364,_T_365};
  assign _T_367 = _T_119_0_bits_data[31];
  assign _T_368 = _T_126_0_data[31];
  assign _T_369 = {_T_367,_T_368};
  assign _T_370 = _T_119_0_lut >> _T_276;
  assign _T_371 = _T_370[0];
  assign _T_372 = _T_119_0_lut >> _T_279;
  assign _T_373 = _T_372[0];
  assign _T_374 = _T_119_0_lut >> _T_282;
  assign _T_375 = _T_374[0];
  assign _T_376 = _T_119_0_lut >> _T_285;
  assign _T_377 = _T_376[0];
  assign _T_378 = _T_119_0_lut >> _T_288;
  assign _T_379 = _T_378[0];
  assign _T_380 = _T_119_0_lut >> _T_291;
  assign _T_381 = _T_380[0];
  assign _T_382 = _T_119_0_lut >> _T_294;
  assign _T_383 = _T_382[0];
  assign _T_384 = _T_119_0_lut >> _T_297;
  assign _T_385 = _T_384[0];
  assign _T_386 = _T_119_0_lut >> _T_300;
  assign _T_387 = _T_386[0];
  assign _T_388 = _T_119_0_lut >> _T_303;
  assign _T_389 = _T_388[0];
  assign _T_390 = _T_119_0_lut >> _T_306;
  assign _T_391 = _T_390[0];
  assign _T_392 = _T_119_0_lut >> _T_309;
  assign _T_393 = _T_392[0];
  assign _T_394 = _T_119_0_lut >> _T_312;
  assign _T_395 = _T_394[0];
  assign _T_396 = _T_119_0_lut >> _T_315;
  assign _T_397 = _T_396[0];
  assign _T_398 = _T_119_0_lut >> _T_318;
  assign _T_399 = _T_398[0];
  assign _T_400 = _T_119_0_lut >> _T_321;
  assign _T_401 = _T_400[0];
  assign _T_402 = _T_119_0_lut >> _T_324;
  assign _T_403 = _T_402[0];
  assign _T_404 = _T_119_0_lut >> _T_327;
  assign _T_405 = _T_404[0];
  assign _T_406 = _T_119_0_lut >> _T_330;
  assign _T_407 = _T_406[0];
  assign _T_408 = _T_119_0_lut >> _T_333;
  assign _T_409 = _T_408[0];
  assign _T_410 = _T_119_0_lut >> _T_336;
  assign _T_411 = _T_410[0];
  assign _T_412 = _T_119_0_lut >> _T_339;
  assign _T_413 = _T_412[0];
  assign _T_414 = _T_119_0_lut >> _T_342;
  assign _T_415 = _T_414[0];
  assign _T_416 = _T_119_0_lut >> _T_345;
  assign _T_417 = _T_416[0];
  assign _T_418 = _T_119_0_lut >> _T_348;
  assign _T_419 = _T_418[0];
  assign _T_420 = _T_119_0_lut >> _T_351;
  assign _T_421 = _T_420[0];
  assign _T_422 = _T_119_0_lut >> _T_354;
  assign _T_423 = _T_422[0];
  assign _T_424 = _T_119_0_lut >> _T_357;
  assign _T_425 = _T_424[0];
  assign _T_426 = _T_119_0_lut >> _T_360;
  assign _T_427 = _T_426[0];
  assign _T_428 = _T_119_0_lut >> _T_363;
  assign _T_429 = _T_428[0];
  assign _T_430 = _T_119_0_lut >> _T_366;
  assign _T_431 = _T_430[0];
  assign _T_432 = _T_119_0_lut >> _T_369;
  assign _T_433 = _T_432[0];
  assign _T_434 = {_T_373,_T_371};
  assign _T_435 = {_T_377,_T_375};
  assign _T_436 = {_T_435,_T_434};
  assign _T_437 = {_T_381,_T_379};
  assign _T_438 = {_T_385,_T_383};
  assign _T_439 = {_T_438,_T_437};
  assign _T_440 = {_T_439,_T_436};
  assign _T_441 = {_T_389,_T_387};
  assign _T_442 = {_T_393,_T_391};
  assign _T_443 = {_T_442,_T_441};
  assign _T_444 = {_T_397,_T_395};
  assign _T_445 = {_T_401,_T_399};
  assign _T_446 = {_T_445,_T_444};
  assign _T_447 = {_T_446,_T_443};
  assign _T_448 = {_T_447,_T_440};
  assign _T_449 = {_T_405,_T_403};
  assign _T_450 = {_T_409,_T_407};
  assign _T_451 = {_T_450,_T_449};
  assign _T_452 = {_T_413,_T_411};
  assign _T_453 = {_T_417,_T_415};
  assign _T_454 = {_T_453,_T_452};
  assign _T_455 = {_T_454,_T_451};
  assign _T_456 = {_T_421,_T_419};
  assign _T_457 = {_T_425,_T_423};
  assign _T_458 = {_T_457,_T_456};
  assign _T_459 = {_T_429,_T_427};
  assign _T_460 = {_T_433,_T_431};
  assign _T_461 = {_T_460,_T_459};
  assign _T_462 = {_T_461,_T_458};
  assign _T_463 = {_T_462,_T_455};
  assign _T_464 = {_T_463,_T_448};
  assign _T_465 = _T_119_0_bits_param[1];
  assign _T_466 = _T_119_0_bits_param[0];
  assign _T_467 = _T_119_0_bits_param[2];
  assign _T_468 = ~ _T_119_0_bits_mask;
  assign _T_469 = _T_119_0_bits_mask[3:1];
  assign _GEN_32 = {{1'd0}, _T_469};
  assign _T_470 = _T_468 | _GEN_32;
  assign _T_471 = ~ _T_470;
  assign _T_476 = {_T_319,_T_295};
  assign _T_477 = {_T_367,_T_343};
  assign _T_478 = {_T_477,_T_476};
  assign _T_483 = {_T_320,_T_296};
  assign _T_484 = {_T_368,_T_344};
  assign _T_485 = {_T_484,_T_483};
  assign _T_486 = _T_478 & _T_471;
  assign _GEN_33 = {{1'd0}, _T_486};
  assign _T_487 = _GEN_33 << 1;
  assign _T_488 = _T_487[3:0];
  assign _T_489 = _T_485 & _T_471;
  assign _GEN_34 = {{1'd0}, _T_489};
  assign _T_490 = _GEN_34 << 1;
  assign _T_491 = _T_490[3:0];
  assign _GEN_35 = {{1'd0}, _T_488};
  assign _T_492 = _GEN_35 << 1;
  assign _T_493 = _T_492[3:0];
  assign _T_494 = _T_488 | _T_493;
  assign _GEN_36 = {{2'd0}, _T_494};
  assign _T_495 = _GEN_36 << 2;
  assign _T_496 = _T_495[3:0];
  assign _T_497 = _T_494 | _T_496;
  assign _T_499 = _T_497[0];
  assign _T_500 = _T_497[1];
  assign _T_501 = _T_497[2];
  assign _T_502 = _T_497[3];
  assign _T_506 = _T_499 ? 8'hff : 8'h0;
  assign _T_510 = _T_500 ? 8'hff : 8'h0;
  assign _T_514 = _T_501 ? 8'hff : 8'h0;
  assign _T_518 = _T_502 ? 8'hff : 8'h0;
  assign _T_519 = {_T_510,_T_506};
  assign _T_520 = {_T_518,_T_514};
  assign _T_521 = {_T_520,_T_519};
  assign _GEN_37 = {{1'd0}, _T_491};
  assign _T_522 = _GEN_37 << 1;
  assign _T_523 = _T_522[3:0];
  assign _T_524 = _T_491 | _T_523;
  assign _GEN_38 = {{2'd0}, _T_524};
  assign _T_525 = _GEN_38 << 2;
  assign _T_526 = _T_525[3:0];
  assign _T_527 = _T_524 | _T_526;
  assign _T_529 = _T_527[0];
  assign _T_530 = _T_527[1];
  assign _T_531 = _T_527[2];
  assign _T_532 = _T_527[3];
  assign _T_536 = _T_529 ? 8'hff : 8'h0;
  assign _T_540 = _T_530 ? 8'hff : 8'h0;
  assign _T_544 = _T_531 ? 8'hff : 8'h0;
  assign _T_548 = _T_532 ? 8'hff : 8'h0;
  assign _T_549 = {_T_540,_T_536};
  assign _T_550 = {_T_548,_T_544};
  assign _T_551 = {_T_550,_T_549};
  assign _T_552 = _T_119_0_bits_mask[0];
  assign _T_553 = _T_119_0_bits_mask[1];
  assign _T_554 = _T_119_0_bits_mask[2];
  assign _T_555 = _T_119_0_bits_mask[3];
  assign _T_559 = _T_552 ? 8'hff : 8'h0;
  assign _T_563 = _T_553 ? 8'hff : 8'h0;
  assign _T_567 = _T_554 ? 8'hff : 8'h0;
  assign _T_571 = _T_555 ? 8'hff : 8'h0;
  assign _T_572 = {_T_563,_T_559};
  assign _T_573 = {_T_571,_T_567};
  assign _T_574 = {_T_573,_T_572};
  assign _T_575 = _T_119_0_bits_data & _T_574;
  assign _T_576 = _T_575 | _T_521;
  assign _T_577 = _T_126_0_data & _T_574;
  assign _T_578 = _T_577 | _T_551;
  assign _T_579 = ~ _T_578;
  assign _T_580 = _T_467 ? _T_578 : _T_579;
  assign _T_581 = _T_576 + _T_580;
  assign _T_582 = _T_581[31:0];
  assign _T_583 = _T_576[31];
  assign _T_584 = _T_465 == _T_583;
  assign _T_586 = _T_578[31];
  assign _T_587 = _T_583 == _T_586;
  assign _T_588 = _T_582[31];
  assign _T_590 = _T_588 == 1'h0;
  assign _T_591 = _T_587 ? _T_590 : _T_584;
  assign _T_592 = _T_466 == _T_591;
  assign _T_593 = _T_592 ? _T_119_0_bits_data : _T_126_0_data;
  assign _T_594 = _T_467 ? _T_582 : _T_593;
  assign _T_595 = _T_119_0_bits_opcode[0];
  assign _T_596 = _T_595 ? _T_464 : _T_594;
  assign _T_602 = _T_268 == 1'h0;
  assign _T_603 = _T_202 | _T_130;
  assign _T_604 = _T_602 & _T_603;
  assign _T_605 = _T_821 & _T_604;
  assign _T_606 = io_in_0_a_valid & _T_604;
  assign _T_608 = _T_202 == 1'h0;
  assign _GEN_0 = _T_608 ? 3'h4 : io_in_0_a_bits_opcode;
  assign _GEN_1 = _T_608 ? 3'h0 : io_in_0_a_bits_param;
  assign _T_659 = _T_119_0_bits_size[0];
  assign _T_661 = 2'h1 << _T_659;
  assign _T_664 = _T_661 | 2'h1;
  assign _T_666 = _T_119_0_bits_size >= 3'h2;
  assign _T_668 = _T_664[1];
  assign _T_669 = _T_119_0_bits_address[1];
  assign _T_671 = _T_669 == 1'h0;
  assign _T_673 = _T_668 & _T_671;
  assign _T_674 = _T_666 | _T_673;
  assign _T_676 = _T_668 & _T_669;
  assign _T_677 = _T_666 | _T_676;
  assign _T_678 = _T_664[0];
  assign _T_679 = _T_119_0_bits_address[0];
  assign _T_681 = _T_679 == 1'h0;
  assign _T_682 = _T_671 & _T_681;
  assign _T_683 = _T_678 & _T_682;
  assign _T_684 = _T_674 | _T_683;
  assign _T_685 = _T_671 & _T_679;
  assign _T_686 = _T_678 & _T_685;
  assign _T_687 = _T_674 | _T_686;
  assign _T_688 = _T_669 & _T_681;
  assign _T_689 = _T_678 & _T_688;
  assign _T_690 = _T_677 | _T_689;
  assign _T_691 = _T_669 & _T_679;
  assign _T_692 = _T_678 & _T_691;
  assign _T_693 = _T_677 | _T_692;
  assign _T_694 = {_T_687,_T_684};
  assign _T_695 = {_T_693,_T_690};
  assign _T_696 = {_T_695,_T_694};
  assign _T_700 = 13'h3f << io_in_0_a_bits_size;
  assign _T_701 = _T_700[5:0];
  assign _T_702 = ~ _T_701;
  assign _T_703 = _T_702[5:2];
  assign _T_704 = io_in_0_a_bits_opcode[2];
  assign _T_706 = _T_704 == 1'h0;
  assign _T_708 = _T_706 ? _T_703 : 4'h0;
  assign _T_713 = _T_711 == 4'h0;
  assign _T_714 = _T_713 & io_out_0_a_ready;
  assign _T_715 = {_T_606,_T_131};
  assign _GEN_39 = {{1'd0}, _T_715};
  assign _T_716 = _GEN_39 << 1;
  assign _T_717 = _T_716[1:0];
  assign _T_718 = _T_715 | _T_717;
  assign _GEN_40 = {{1'd0}, _T_718};
  assign _T_720 = _GEN_40 << 1;
  assign _T_721 = _T_720[1:0];
  assign _T_722 = ~ _T_721;
  assign _T_723 = _T_722[0];
  assign _T_724 = _T_722[1];
  assign _T_732 = _T_723 & _T_131;
  assign _T_733 = _T_724 & _T_606;
  assign _T_743 = _T_732 | _T_733;
  assign _T_747 = _T_732 == 1'h0;
  assign _T_752 = _T_733 == 1'h0;
  assign _T_753 = _T_747 | _T_752;
  assign _T_755 = _T_753 | reset;
  assign _T_757 = _T_755 == 1'h0;
  assign _T_758 = _T_131 | _T_606;
  assign _T_760 = _T_758 == 1'h0;
  assign _T_762 = _T_760 | _T_743;
  assign _T_763 = _T_762 | reset;
  assign _T_765 = _T_763 == 1'h0;
  assign _T_769 = _T_733 ? _T_708 : 4'h0;
  assign _T_771 = io_out_0_a_ready & io_out_0_a_valid;
  assign _GEN_41 = {{3'd0}, _T_771};
  assign _T_772 = _T_711 - _GEN_41;
  assign _T_773 = $unsigned(_T_772);
  assign _T_774 = _T_773[3:0];
  assign _T_775 = _T_714 ? _T_769 : _T_774;
  assign _T_804_0 = _T_713 ? _T_732 : _T_793_0;
  assign _T_804_1 = _T_713 ? _T_733 : _T_793_1;
  assign _T_812_0 = _T_713 ? _T_723 : _T_793_0;
  assign _T_812_1 = _T_713 ? _T_724 : _T_793_1;
  assign _T_820 = io_out_0_a_ready & _T_812_0;
  assign _T_821 = io_out_0_a_ready & _T_812_1;
  assign _T_825 = _T_793_0 ? _T_131 : 1'h0;
  assign _T_827 = _T_793_1 ? _T_606 : 1'h0;
  assign _T_828 = _T_825 | _T_827;
  assign _T_831 = _T_713 ? _T_758 : _T_828;
  assign _T_833 = {_T_119_0_bits_address,_T_696};
  assign _T_834 = {_T_833,_T_596};
  assign _T_835 = {_T_119_0_bits_size,_T_119_0_bits_source};
  assign _T_837 = {6'h0,_T_835};
  assign _T_838 = {_T_837,_T_834};
  assign _T_840 = _T_804_0 ? _T_838 : 82'h0;
  assign _T_841 = {io_in_0_a_bits_address,io_in_0_a_bits_mask};
  assign _T_842 = {_T_841,io_in_0_a_bits_data};
  assign _T_843 = {io_in_0_a_bits_size,io_in_0_a_bits_source};
  assign _T_844 = {_GEN_0,_GEN_1};
  assign _T_845 = {_T_844,_T_843};
  assign _T_846 = {_T_845,_T_842};
  assign _T_848 = _T_804_1 ? _T_846 : 82'h0;
  assign _T_849 = _T_840 | _T_848;
  assign _T_854 = _T_849[31:0];
  assign _T_855 = _T_849[35:32];
  assign _T_856 = _T_849[67:36];
  assign _T_857 = _T_849[72:68];
  assign _T_858 = _T_849[75:73];
  assign _T_859 = _T_849[78:76];
  assign _T_860 = _T_849[81:79];
  assign _T_861 = _T_821 & _T_606;
  assign _T_864 = _T_861 & _T_608;
  assign _T_865 = io_in_0_a_bits_param[1:0];
  assign _GEN_42 = {{1'd0}, _T_865};
  assign _T_875 = 3'h3 == _GEN_42;
  assign _T_876 = _T_875 ? 4'hc : 4'h0;
  assign _T_877 = 3'h0 == _GEN_42;
  assign _T_878 = _T_877 ? 4'h6 : _T_876;
  assign _T_879 = 3'h1 == _GEN_42;
  assign _T_880 = _T_879 ? 4'he : _T_878;
  assign _T_881 = 3'h2 == _GEN_42;
  assign _T_882 = _T_881 ? 4'h8 : _T_880;
  assign _GEN_2 = _T_130 ? _T_263 : _T_119_0_fifoId;
  assign _GEN_3 = _T_130 ? io_in_0_a_bits_opcode : _T_119_0_bits_opcode;
  assign _GEN_4 = _T_130 ? io_in_0_a_bits_param : _T_119_0_bits_param;
  assign _GEN_5 = _T_130 ? io_in_0_a_bits_size : _T_119_0_bits_size;
  assign _GEN_6 = _T_130 ? io_in_0_a_bits_source : _T_119_0_bits_source;
  assign _GEN_7 = _T_130 ? io_in_0_a_bits_address : _T_119_0_bits_address;
  assign _GEN_8 = _T_130 ? io_in_0_a_bits_mask : _T_119_0_bits_mask;
  assign _GEN_9 = _T_130 ? io_in_0_a_bits_data : _T_119_0_bits_data;
  assign _GEN_10 = _T_130 ? _T_882 : _T_119_0_lut;
  assign _GEN_11 = _T_130 ? 2'h3 : _T_108_0_state;
  assign _GEN_12 = _T_864 ? _GEN_2 : _T_119_0_fifoId;
  assign _GEN_13 = _T_864 ? _GEN_3 : _T_119_0_bits_opcode;
  assign _GEN_14 = _T_864 ? _GEN_4 : _T_119_0_bits_param;
  assign _GEN_15 = _T_864 ? _GEN_5 : _T_119_0_bits_size;
  assign _GEN_16 = _T_864 ? _GEN_6 : _T_119_0_bits_source;
  assign _GEN_17 = _T_864 ? _GEN_7 : _T_119_0_bits_address;
  assign _GEN_18 = _T_864 ? _GEN_8 : _T_119_0_bits_mask;
  assign _GEN_19 = _T_864 ? _GEN_9 : _T_119_0_bits_data;
  assign _GEN_20 = _T_864 ? _GEN_10 : _T_119_0_lut;
  assign _GEN_21 = _T_864 ? _GEN_11 : _T_108_0_state;
  assign _T_883 = _T_820 & _T_131;
  assign _GEN_22 = _T_131 ? 2'h1 : _GEN_21;
  assign _GEN_23 = _T_883 ? _GEN_22 : _GEN_21;
  assign _T_884 = io_out_0_d_ready & io_out_0_d_valid;
  assign _T_887 = 13'h3f << io_out_0_d_bits_size;
  assign _T_888 = _T_887[5:0];
  assign _T_889 = ~ _T_888;
  assign _T_890 = _T_889[5:2];
  assign _T_891 = io_out_0_d_bits_opcode[0];
  assign _T_893 = _T_891 ? _T_890 : 4'h0;
  assign _T_898 = _T_896 - 4'h1;
  assign _T_899 = $unsigned(_T_898);
  assign _T_900 = _T_899[3:0];
  assign _T_902 = _T_896 == 4'h0;
  assign _T_911 = _T_902 ? _T_893 : _T_900;
  assign _GEN_24 = _T_884 ? _T_911 : _T_896;
  assign _T_912 = _T_119_0_bits_source == io_in_0_d_bits_source;
  assign _T_913 = _T_912 & _T_135;
  assign _T_918 = io_out_0_d_bits_opcode == 3'h1;
  assign _T_920 = io_out_0_d_bits_opcode == 3'h0;
  assign _T_922 = _T_884 & _T_902;
  assign _T_923 = _T_913 & _T_918;
  assign _GEN_25 = _T_923 ? io_out_0_d_bits_data : _T_126_0_data;
  assign _T_924 = _T_918 ? 2'h2 : 2'h0;
  assign _GEN_26 = _T_913 ? _T_924 : _GEN_23;
  assign _GEN_27 = _T_922 ? _GEN_25 : _T_126_0_data;
  assign _GEN_28 = _T_922 ? _GEN_26 : _GEN_23;
  assign _T_925 = _T_902 & _T_918;
  assign _T_926 = _T_925 & _T_913;
  assign _T_927 = _T_902 & _T_920;
  assign _T_928 = _T_927 & _T_913;
  assign _T_930 = _T_926 == 1'h0;
  assign _T_931 = io_out_0_d_valid & _T_930;
  assign _T_932 = io_in_0_d_ready | _T_926;
  assign _GEN_29 = _T_928 ? 3'h1 : io_out_0_d_bits_opcode;
  assign _GEN_30 = _T_928 ? _T_126_0_data : io_out_0_d_bits_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_108_0_state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_119_0_bits_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_119_0_bits_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_119_0_bits_size = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_119_0_bits_source = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_119_0_bits_address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_119_0_bits_mask = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_119_0_bits_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_119_0_fifoId = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_119_0_lut = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_126_0_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_711 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_793_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_793_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_896 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_108_0_state <= 2'h0;
    end else begin
      if (_T_922) begin
        if (_T_913) begin
          if (_T_918) begin
            _T_108_0_state <= 2'h2;
          end else begin
            _T_108_0_state <= 2'h0;
          end
        end else begin
          if (_T_883) begin
            if (_T_131) begin
              _T_108_0_state <= 2'h1;
            end else begin
              if (_T_864) begin
                if (_T_130) begin
                  _T_108_0_state <= 2'h3;
                end
              end
            end
          end else begin
            if (_T_864) begin
              if (_T_130) begin
                _T_108_0_state <= 2'h3;
              end
            end
          end
        end
      end else begin
        if (_T_883) begin
          if (_T_131) begin
            _T_108_0_state <= 2'h1;
          end else begin
            if (_T_864) begin
              if (_T_130) begin
                _T_108_0_state <= 2'h3;
              end
            end
          end
        end else begin
          if (_T_864) begin
            if (_T_130) begin
              _T_108_0_state <= 2'h3;
            end
          end
        end
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_opcode <= io_in_0_a_bits_opcode;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_param <= io_in_0_a_bits_param;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_size <= io_in_0_a_bits_size;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_source <= io_in_0_a_bits_source;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_address <= io_in_0_a_bits_address;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_mask <= io_in_0_a_bits_mask;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_bits_data <= io_in_0_a_bits_data;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        _T_119_0_fifoId <= _T_263;
      end
    end
    if (_T_864) begin
      if (_T_130) begin
        if (_T_881) begin
          _T_119_0_lut <= 4'h8;
        end else begin
          if (_T_879) begin
            _T_119_0_lut <= 4'he;
          end else begin
            if (_T_877) begin
              _T_119_0_lut <= 4'h6;
            end else begin
              if (_T_875) begin
                _T_119_0_lut <= 4'hc;
              end else begin
                _T_119_0_lut <= 4'h0;
              end
            end
          end
        end
      end
    end
    if (_T_922) begin
      if (_T_923) begin
        _T_126_0_data <= io_out_0_d_bits_data;
      end
    end
    if (reset) begin
      _T_711 <= 4'h0;
    end else begin
      if (_T_714) begin
        if (_T_733) begin
          if (_T_706) begin
            _T_711 <= _T_703;
          end else begin
            _T_711 <= 4'h0;
          end
        end else begin
          _T_711 <= 4'h0;
        end
      end else begin
        _T_711 <= _T_774;
      end
    end
    if (reset) begin
      _T_793_0 <= 1'h0;
    end else begin
      if (_T_713) begin
        _T_793_0 <= _T_732;
      end
    end
    if (reset) begin
      _T_793_1 <= 1'h0;
    end else begin
      if (_T_713) begin
        _T_793_1 <= _T_733;
      end
    end
    if (reset) begin
      _T_896 <= 4'h0;
    end else begin
      if (_T_884) begin
        if (_T_902) begin
          if (_T_891) begin
            _T_896 <= _T_890;
          end else begin
            _T_896 <= 4'h0;
          end
        end else begin
          _T_896 <= _T_900;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_757) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_757) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_765) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_765) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LevelGateway(
  input   clock,
  input   reset,
  input   io_interrupt,
  output  io_plic_valid,
  input   io_plic_ready,
  input   io_plic_complete
);
  reg  inFlight;
  reg [31:0] _RAND_0;
  wire  _T_8;
  wire  _GEN_0;
  wire  _GEN_1;
  wire  _T_12;
  wire  _T_13;
  assign io_plic_valid = _T_13;
  assign _T_8 = io_interrupt & io_plic_ready;
  assign _GEN_0 = _T_8 ? 1'h1 : inFlight;
  assign _GEN_1 = io_plic_complete ? 1'h0 : _GEN_0;
  assign _T_12 = inFlight == 1'h0;
  assign _T_13 = io_interrupt & _T_12;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  inFlight = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      inFlight <= 1'h0;
    end else begin
      if (io_plic_complete) begin
        inFlight <= 1'h0;
      end else begin
        if (_T_8) begin
          inFlight <= 1'h1;
        end
      end
    end
  end
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_read,
  input  [23:0] io_enq_bits_index,
  input  [31:0] io_enq_bits_data,
  input  [3:0]  io_enq_bits_mask,
  input  [11:0] io_enq_bits_extra,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_read,
  output [23:0] io_deq_bits_index,
  output [31:0] io_deq_bits_data,
  output [3:0]  io_deq_bits_mask,
  output [11:0] io_deq_bits_extra
);
  reg  ram_read [0:0];
  reg [31:0] _RAND_0;
  wire  ram_read__T_35_data;
  wire  ram_read__T_35_addr;
  wire  ram_read__T_26_data;
  wire  ram_read__T_26_addr;
  wire  ram_read__T_26_mask;
  wire  ram_read__T_26_en;
  reg [23:0] ram_index [0:0];
  reg [31:0] _RAND_1;
  wire [23:0] ram_index__T_35_data;
  wire  ram_index__T_35_addr;
  wire [23:0] ram_index__T_26_data;
  wire  ram_index__T_26_addr;
  wire  ram_index__T_26_mask;
  wire  ram_index__T_26_en;
  reg [31:0] ram_data [0:0];
  reg [31:0] _RAND_2;
  wire [31:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [31:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg [3:0] ram_mask [0:0];
  reg [31:0] _RAND_3;
  wire [3:0] ram_mask__T_35_data;
  wire  ram_mask__T_35_addr;
  wire [3:0] ram_mask__T_26_data;
  wire  ram_mask__T_26_addr;
  wire  ram_mask__T_26_mask;
  wire  ram_mask__T_26_en;
  reg [11:0] ram_extra [0:0];
  reg [31:0] _RAND_4;
  wire [11:0] ram_extra__T_35_data;
  wire  ram_extra__T_35_addr;
  wire [11:0] ram_extra__T_26_data;
  wire  ram_extra__T_26_addr;
  wire  ram_extra__T_26_mask;
  wire  ram_extra__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_8;
  wire  _T_31;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _T_31;
  assign io_deq_bits_read = ram_read__T_35_data;
  assign io_deq_bits_index = ram_index__T_35_data;
  assign io_deq_bits_data = ram_data__T_35_data;
  assign io_deq_bits_mask = ram_mask__T_35_data;
  assign io_deq_bits_extra = ram_extra__T_35_data;
  assign ram_read__T_35_addr = 1'h0;
  assign ram_read__T_35_data = ram_read[ram_read__T_35_addr];
  assign ram_read__T_26_data = io_enq_bits_read;
  assign ram_read__T_26_addr = 1'h0;
  assign ram_read__T_26_mask = _T_21;
  assign ram_read__T_26_en = _T_21;
  assign ram_index__T_35_addr = 1'h0;
  assign ram_index__T_35_data = ram_index[ram_index__T_35_addr];
  assign ram_index__T_26_data = io_enq_bits_index;
  assign ram_index__T_26_addr = 1'h0;
  assign ram_index__T_26_mask = _T_21;
  assign ram_index__T_26_en = _T_21;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _T_21;
  assign ram_data__T_26_en = _T_21;
  assign ram_mask__T_35_addr = 1'h0;
  assign ram_mask__T_35_data = ram_mask[ram_mask__T_35_addr];
  assign ram_mask__T_26_data = io_enq_bits_mask;
  assign ram_mask__T_26_addr = 1'h0;
  assign ram_mask__T_26_mask = _T_21;
  assign ram_mask__T_26_en = _T_21;
  assign ram_extra__T_35_addr = 1'h0;
  assign ram_extra__T_35_data = ram_extra[ram_extra__T_35_addr];
  assign ram_extra__T_26_data = io_enq_bits_extra;
  assign ram_extra__T_26_addr = 1'h0;
  assign ram_extra__T_26_mask = _T_21;
  assign ram_extra__T_26_en = _T_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _T_21 != _T_23;
  assign _GEN_8 = _T_29 ? _T_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_read[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_index[initvar] = _RAND_1[23:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_mask[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_extra[initvar] = _RAND_4[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_read__T_26_en & ram_read__T_26_mask) begin
      ram_read[ram_read__T_26_addr] <= ram_read__T_26_data;
    end
    if(ram_index__T_26_en & ram_index__T_26_mask) begin
      ram_index[ram_index__T_26_addr] <= ram_index__T_26_data;
    end
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if(ram_mask__T_26_en & ram_mask__T_26_mask) begin
      ram_mask[ram_mask__T_26_addr] <= ram_mask__T_26_data;
    end
    if(ram_extra__T_26_en & ram_extra__T_26_mask) begin
      ram_extra[ram_extra__T_26_addr] <= ram_extra__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        maybe_full <= _T_21;
      end
    end
  end
endmodule
module TLPLIC_plic(
  input         clock,
  input         reset,
  output        io_tl_in_0_a_ready,
  input         io_tl_in_0_a_valid,
  input  [2:0]  io_tl_in_0_a_bits_opcode,
  input  [1:0]  io_tl_in_0_a_bits_size,
  input  [9:0]  io_tl_in_0_a_bits_source,
  input  [27:0] io_tl_in_0_a_bits_address,
  input  [3:0]  io_tl_in_0_a_bits_mask,
  input  [31:0] io_tl_in_0_a_bits_data,
  input         io_tl_in_0_d_ready,
  output        io_tl_in_0_d_valid,
  output [2:0]  io_tl_in_0_d_bits_opcode,
  output [1:0]  io_tl_in_0_d_bits_param,
  output [1:0]  io_tl_in_0_d_bits_size,
  output [9:0]  io_tl_in_0_d_bits_source,
  output        io_tl_in_0_d_bits_sink,
  output [31:0] io_tl_in_0_d_bits_data,
  output        io_tl_in_0_d_bits_error,
  input         io_devices_0_0,
  input         io_devices_0_1,
  output        io_harts_0_0
);
  wire  LevelGateway_clock;
  wire  LevelGateway_reset;
  wire  LevelGateway_io_interrupt;
  wire  LevelGateway_io_plic_valid;
  wire  LevelGateway_io_plic_ready;
  wire  LevelGateway_io_plic_complete;
  wire  LevelGateway_1_clock;
  wire  LevelGateway_1_reset;
  wire  LevelGateway_1_io_interrupt;
  wire  LevelGateway_1_io_plic_valid;
  wire  LevelGateway_1_io_plic_ready;
  wire  LevelGateway_1_io_plic_complete;
  wire  LevelGateway_2_clock;
  wire  LevelGateway_2_reset;
  wire  LevelGateway_2_io_interrupt;
  wire  LevelGateway_2_io_plic_valid;
  wire  LevelGateway_2_io_plic_ready;
  wire  LevelGateway_2_io_plic_complete;
  wire  gateways_1_valid;
  wire  gateways_2_valid;
  reg [1:0] priority_0;
  reg [31:0] _RAND_0;
  reg [1:0] priority_1;
  reg [31:0] _RAND_1;
  reg [1:0] priority_2;
  reg [31:0] _RAND_2;
  reg [1:0] threshold_0;
  reg [31:0] _RAND_3;
  reg  pending_0;
  reg [31:0] _RAND_4;
  reg  pending_1;
  reg [31:0] _RAND_5;
  reg  pending_2;
  reg [31:0] _RAND_6;
  reg  enables_0_0;
  reg [31:0] _RAND_7;
  reg  enables_0_1;
  reg [31:0] _RAND_8;
  reg  enables_0_2;
  reg [31:0] _RAND_9;
  reg [1:0] maxDevs_0;
  reg [31:0] _RAND_10;
  wire  _T_219;
  wire [2:0] _T_220;
  wire  _T_221;
  wire [2:0] _T_222;
  wire  _T_225;
  wire [2:0] _T_228;
  wire  _T_229;
  wire  _T_231;
  wire [2:0] _T_234;
  wire [1:0] _T_235;
  reg [2:0] _T_237;
  reg [31:0] _RAND_11;
  wire [2:0] _T_239;
  wire  _T_240;
  wire [1:0] _T_248;
  wire [1:0] _T_249;
  wire  _T_250;
  wire  _T_251;
  wire  _T_253;
  wire  _T_254;
  wire  _T_256;
  wire [3:0] _T_259;
  wire [2:0] _T_260;
  wire [2:0] _T_262;
  wire  _T_269;
  wire  _T_270;
  wire  _T_279;
  wire  _T_284;
  wire  _T_285;
  wire  _T_287;
  wire  _GEN_8;
  wire  _T_289;
  wire  _T_290;
  wire  _T_292;
  wire  _GEN_9;
  wire [1:0] _T_300;
  wire [1:0] _T_301;
  wire  _T_302;
  wire  _T_303;
  wire  _T_305;
  wire  _T_306;
  wire  _T_308;
  wire [3:0] _T_312;
  wire [2:0] _T_313;
  wire [2:0] completedDevs;
  wire  _T_315;
  wire  _T_316;
  wire  _T_317;
  wire [23:0] _T_323_bits_index;
  wire  _T_328;
  wire [25:0] _T_329;
  wire [11:0] _T_330;
  wire  _T_336_bits_read;
  wire [11:0] _T_336_bits_extra;
  wire  _T_345_ready;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire  Queue_io_enq_bits_read;
  wire [23:0] Queue_io_enq_bits_index;
  wire [31:0] Queue_io_enq_bits_data;
  wire [3:0] Queue_io_enq_bits_mask;
  wire [11:0] Queue_io_enq_bits_extra;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire  Queue_io_deq_bits_read;
  wire [23:0] Queue_io_deq_bits_index;
  wire [31:0] Queue_io_deq_bits_data;
  wire [3:0] Queue_io_deq_bits_mask;
  wire [11:0] Queue_io_deq_bits_extra;
  wire [23:0] _T_421;
  wire [23:0] _T_422;
  wire  _T_424;
  wire [23:0] _T_430;
  wire [23:0] _T_431;
  wire  _T_433;
  wire [23:0] _T_439;
  wire [23:0] _T_440;
  wire  _T_442;
  wire [23:0] _T_448;
  wire [23:0] _T_449;
  wire  _T_451;
  wire [23:0] _T_457;
  wire [23:0] _T_458;
  wire  _T_460;
  wire [23:0] _T_466;
  wire [23:0] _T_467;
  wire  _T_469;
  wire [23:0] _T_475;
  wire [23:0] _T_476;
  wire  _T_478;
  wire  _T_602;
  wire  _T_603;
  wire  _T_604;
  wire  _T_605;
  wire [7:0] _T_609;
  wire [7:0] _T_613;
  wire [7:0] _T_617;
  wire [7:0] _T_621;
  wire [15:0] _T_622;
  wire [15:0] _T_623;
  wire [31:0] _T_624;
  wire  _T_672;
  wire  _T_676;
  wire  _T_678;
  wire  _T_685;
  wire [1:0] _GEN_205;
  wire [1:0] _T_700;
  wire [1:0] _GEN_206;
  wire [1:0] _T_704;
  wire  _T_712;
  wire  _T_716;
  wire  _T_718;
  wire  _T_725;
  wire [2:0] _GEN_207;
  wire [2:0] _T_740;
  wire [2:0] _GEN_208;
  wire [2:0] _T_744;
  wire  _T_754;
  wire [31:0] _T_756;
  wire  _T_758;
  wire [31:0] _T_765;
  wire [31:0] _T_783;
  wire  _T_800;
  wire  _T_804;
  wire [1:0] _T_807;
  wire  _T_808;
  wire  _T_809;
  wire  _T_811;
  wire [1:0] _T_812;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _T_815;
  wire [31:0] _T_832;
  wire  _T_853;
  wire [31:0] _GEN_13;
  wire [31:0] _T_872;
  wire  _T_893;
  wire [31:0] _GEN_14;
  wire [31:0] _T_912;
  wire  _T_933;
  wire [31:0] _GEN_15;
  wire [31:0] _T_952;
  wire  _T_1013;
  wire  _GEN_17;
  wire [1:0] _GEN_209;
  wire [1:0] _T_1029;
  wire [1:0] _GEN_210;
  wire [1:0] _T_1033;
  wire  _T_1053;
  wire  _GEN_18;
  wire [2:0] _GEN_211;
  wire [2:0] _T_1069;
  wire [2:0] _GEN_212;
  wire [2:0] _T_1073;
  wire  _T_1102;
  wire  _T_1103;
  wire  _T_1112;
  wire  _T_1113;
  wire  _T_1121;
  wire [1:0] _T_1126;
  wire [1:0] _T_1127;
  wire [2:0] _T_1128;
  wire [4:0] _T_1129;
  wire [31:0] _T_1165;
  wire  _T_1167;
  wire  _T_1168;
  wire  _T_1174;
  wire  _T_1182;
  wire  _T_1183;
  wire  _T_1790;
  wire  _T_1791;
  wire  _T_1930;
  wire  _T_1931;
  wire  _T_2087;
  wire  _T_2088;
  wire  _T_2099;
  wire  _T_2100;
  wire  _T_2107;
  wire  _T_2108;
  wire  _T_2155;
  wire  _T_2156;
  wire  _T_2219;
  wire  _T_2220;
  wire  _T_2227;
  wire  _T_2228;
  wire  _T_2391;
  wire [31:0] _T_2432_4;
  wire [31:0] _T_2432_8;
  wire  _GEN_143;
  wire  _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire  _GEN_147;
  wire  _GEN_148;
  wire  _GEN_149;
  wire  _GEN_150;
  wire  _GEN_151;
  wire  _GEN_152;
  wire  _GEN_153;
  wire  _GEN_154;
  wire  _GEN_155;
  wire  _GEN_156;
  wire  _GEN_157;
  wire  _GEN_158;
  wire  _GEN_159;
  wire  _GEN_160;
  wire  _GEN_161;
  wire  _GEN_162;
  wire  _GEN_163;
  wire  _GEN_164;
  wire  _GEN_165;
  wire  _GEN_166;
  wire  _GEN_167;
  wire  _GEN_168;
  wire  _GEN_169;
  wire  _GEN_170;
  wire  _GEN_171;
  wire  _GEN_172;
  wire  _GEN_173;
  wire [31:0] _GEN_174;
  wire [31:0] _GEN_175;
  wire [31:0] _GEN_176;
  wire [31:0] _GEN_177;
  wire [31:0] _GEN_178;
  wire [31:0] _GEN_179;
  wire [31:0] _GEN_180;
  wire [31:0] _GEN_181;
  wire [31:0] _GEN_182;
  wire [31:0] _GEN_183;
  wire [31:0] _GEN_184;
  wire [31:0] _GEN_185;
  wire [31:0] _GEN_186;
  wire [31:0] _GEN_187;
  wire [31:0] _GEN_188;
  wire [31:0] _GEN_189;
  wire [31:0] _GEN_190;
  wire [31:0] _GEN_191;
  wire [31:0] _GEN_192;
  wire [31:0] _GEN_193;
  wire [31:0] _GEN_194;
  wire [31:0] _GEN_195;
  wire [31:0] _GEN_196;
  wire [31:0] _GEN_197;
  wire [31:0] _GEN_198;
  wire [31:0] _GEN_199;
  wire [31:0] _GEN_200;
  wire [31:0] _GEN_201;
  wire [31:0] _GEN_202;
  wire [31:0] _GEN_203;
  wire [31:0] _GEN_204;
  wire [31:0] _T_2469;
  wire [9:0] _T_2470;
  wire [1:0] _T_2471;
  LevelGateway LevelGateway (
    .clock(LevelGateway_clock),
    .reset(LevelGateway_reset),
    .io_interrupt(LevelGateway_io_interrupt),
    .io_plic_valid(LevelGateway_io_plic_valid),
    .io_plic_ready(LevelGateway_io_plic_ready),
    .io_plic_complete(LevelGateway_io_plic_complete)
  );
  LevelGateway LevelGateway_1 (
    .clock(LevelGateway_1_clock),
    .reset(LevelGateway_1_reset),
    .io_interrupt(LevelGateway_1_io_interrupt),
    .io_plic_valid(LevelGateway_1_io_plic_valid),
    .io_plic_ready(LevelGateway_1_io_plic_ready),
    .io_plic_complete(LevelGateway_1_io_plic_complete)
  );
  LevelGateway LevelGateway_2 (
    .clock(LevelGateway_2_clock),
    .reset(LevelGateway_2_reset),
    .io_interrupt(LevelGateway_2_io_interrupt),
    .io_plic_valid(LevelGateway_2_io_plic_valid),
    .io_plic_ready(LevelGateway_2_io_plic_ready),
    .io_plic_complete(LevelGateway_2_io_plic_complete)
  );
  Queue_8 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_read(Queue_io_enq_bits_read),
    .io_enq_bits_index(Queue_io_enq_bits_index),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_extra(Queue_io_enq_bits_extra),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_read(Queue_io_deq_bits_read),
    .io_deq_bits_index(Queue_io_deq_bits_index),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_extra(Queue_io_deq_bits_extra)
  );
  assign io_tl_in_0_a_ready = _T_345_ready;
  assign io_tl_in_0_d_valid = _T_2391;
  assign io_tl_in_0_d_bits_opcode = {{2'd0}, _T_336_bits_read};
  assign io_tl_in_0_d_bits_param = 2'h0;
  assign io_tl_in_0_d_bits_size = _T_2471;
  assign io_tl_in_0_d_bits_source = _T_2470;
  assign io_tl_in_0_d_bits_sink = 1'h0;
  assign io_tl_in_0_d_bits_data = _T_2469;
  assign io_tl_in_0_d_bits_error = 1'h0;
  assign io_harts_0_0 = _T_240;
  assign LevelGateway_clock = clock;
  assign LevelGateway_reset = reset;
  assign LevelGateway_io_interrupt = 1'h0;
  assign LevelGateway_io_plic_ready = _T_279;
  assign LevelGateway_io_plic_complete = _T_315;
  assign LevelGateway_1_clock = clock;
  assign LevelGateway_1_reset = reset;
  assign LevelGateway_1_io_interrupt = io_devices_0_0;
  assign LevelGateway_1_io_plic_ready = _T_284;
  assign LevelGateway_1_io_plic_complete = _T_316;
  assign LevelGateway_2_clock = clock;
  assign LevelGateway_2_reset = reset;
  assign LevelGateway_2_io_interrupt = io_devices_0_1;
  assign LevelGateway_2_io_plic_ready = _T_289;
  assign LevelGateway_2_io_plic_complete = _T_317;
  assign gateways_1_valid = LevelGateway_1_io_plic_valid;
  assign gateways_2_valid = LevelGateway_2_io_plic_valid;
  assign _T_219 = pending_1 & enables_0_1;
  assign _T_220 = {_T_219,priority_1};
  assign _T_221 = pending_2 & enables_0_2;
  assign _T_222 = {_T_221,priority_2};
  assign _T_225 = 3'h4 >= _T_220;
  assign _T_228 = _T_225 ? 3'h4 : _T_220;
  assign _T_229 = _T_225 ? 1'h0 : 1'h1;
  assign _T_231 = _T_228 >= _T_222;
  assign _T_234 = _T_231 ? _T_228 : _T_222;
  assign _T_235 = _T_231 ? {{1'd0}, _T_229} : 2'h2;
  assign _T_239 = {1'h1,threshold_0};
  assign _T_240 = _T_237 > _T_239;
  assign _T_248 = _T_800 - 1'h1;
  assign _T_249 = $unsigned(_T_248);
  assign _T_250 = _T_249[0:0];
  assign _T_251 = _T_800 & _T_250;
  assign _T_253 = _T_251 == 1'h0;
  assign _T_254 = _T_253 | reset;
  assign _T_256 = _T_254 == 1'h0;
  assign _T_259 = 4'h1 << maxDevs_0;
  assign _T_260 = _T_259[2:0];
  assign _T_262 = _T_800 ? _T_260 : 3'h0;
  assign _T_269 = _T_262[1];
  assign _T_270 = _T_262[2];
  assign _T_279 = pending_0 == 1'h0;
  assign _T_284 = pending_1 == 1'h0;
  assign _T_285 = _T_269 | gateways_1_valid;
  assign _T_287 = _T_269 == 1'h0;
  assign _GEN_8 = _T_285 ? _T_287 : pending_1;
  assign _T_289 = pending_2 == 1'h0;
  assign _T_290 = _T_270 | gateways_2_valid;
  assign _T_292 = _T_270 == 1'h0;
  assign _GEN_9 = _T_290 ? _T_292 : pending_2;
  assign _T_300 = _T_815 - 1'h1;
  assign _T_301 = $unsigned(_T_300);
  assign _T_302 = _T_301[0:0];
  assign _T_303 = _T_815 & _T_302;
  assign _T_305 = _T_303 == 1'h0;
  assign _T_306 = _T_305 | reset;
  assign _T_308 = _T_306 == 1'h0;
  assign _T_312 = 4'h1 << _T_812;
  assign _T_313 = _T_312[2:0];
  assign completedDevs = _T_815 ? _T_313 : 3'h0;
  assign _T_315 = completedDevs[0];
  assign _T_316 = completedDevs[1];
  assign _T_317 = completedDevs[2];
  assign _T_323_bits_index = _T_329[23:0];
  assign _T_328 = io_tl_in_0_a_bits_opcode == 3'h4;
  assign _T_329 = io_tl_in_0_a_bits_address[27:2];
  assign _T_330 = {io_tl_in_0_a_bits_source,io_tl_in_0_a_bits_size};
  assign _T_336_bits_read = Queue_io_deq_bits_read;
  assign _T_336_bits_extra = Queue_io_deq_bits_extra;
  assign _T_345_ready = Queue_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_tl_in_0_a_valid;
  assign Queue_io_enq_bits_read = _T_328;
  assign Queue_io_enq_bits_index = _T_323_bits_index;
  assign Queue_io_enq_bits_data = io_tl_in_0_a_bits_data;
  assign Queue_io_enq_bits_mask = io_tl_in_0_a_bits_mask;
  assign Queue_io_enq_bits_extra = _T_330;
  assign Queue_io_deq_ready = io_tl_in_0_d_ready;
  assign _T_421 = Queue_io_deq_bits_index ^ 24'h400;
  assign _T_422 = _T_421 & 24'hf7f3fc;
  assign _T_424 = _T_422 == 24'h0;
  assign _T_430 = Queue_io_deq_bits_index;
  assign _T_431 = _T_430 & 24'hf7f3fc;
  assign _T_433 = _T_431 == 24'h0;
  assign _T_439 = Queue_io_deq_bits_index ^ 24'h80001;
  assign _T_440 = _T_439 & 24'hf7f3fc;
  assign _T_442 = _T_440 == 24'h0;
  assign _T_448 = Queue_io_deq_bits_index ^ 24'h1;
  assign _T_449 = _T_448 & 24'hf7f3fc;
  assign _T_451 = _T_449 == 24'h0;
  assign _T_457 = Queue_io_deq_bits_index ^ 24'h2;
  assign _T_458 = _T_457 & 24'hf7f3fc;
  assign _T_460 = _T_458 == 24'h0;
  assign _T_466 = Queue_io_deq_bits_index ^ 24'h80000;
  assign _T_467 = _T_466 & 24'hf7f3fc;
  assign _T_469 = _T_467 == 24'h0;
  assign _T_475 = Queue_io_deq_bits_index ^ 24'h800;
  assign _T_476 = _T_475 & 24'hf7f3fc;
  assign _T_478 = _T_476 == 24'h0;
  assign _T_602 = Queue_io_deq_bits_mask[0];
  assign _T_603 = Queue_io_deq_bits_mask[1];
  assign _T_604 = Queue_io_deq_bits_mask[2];
  assign _T_605 = Queue_io_deq_bits_mask[3];
  assign _T_609 = _T_602 ? 8'hff : 8'h0;
  assign _T_613 = _T_603 ? 8'hff : 8'h0;
  assign _T_617 = _T_604 ? 8'hff : 8'h0;
  assign _T_621 = _T_605 ? 8'hff : 8'h0;
  assign _T_622 = {_T_613,_T_609};
  assign _T_623 = {_T_621,_T_617};
  assign _T_624 = {_T_623,_T_622};
  assign _T_672 = _T_624[1];
  assign _T_676 = ~ _T_672;
  assign _T_678 = _T_676 == 1'h0;
  assign _T_685 = Queue_io_deq_bits_data[1];
  assign _GEN_205 = {{1'd0}, pending_1};
  assign _T_700 = _GEN_205 << 1;
  assign _GEN_206 = {{1'd0}, pending_0};
  assign _T_704 = _GEN_206 | _T_700;
  assign _T_712 = _T_624[2];
  assign _T_716 = ~ _T_712;
  assign _T_718 = _T_716 == 1'h0;
  assign _T_725 = Queue_io_deq_bits_data[2];
  assign _GEN_207 = {{2'd0}, pending_2};
  assign _T_740 = _GEN_207 << 2;
  assign _GEN_208 = {{1'd0}, _T_704};
  assign _T_744 = _GEN_208 | _T_740;
  assign _T_754 = _T_624 != 32'h0;
  assign _T_756 = ~ _T_624;
  assign _T_758 = _T_756 == 32'h0;
  assign _T_765 = Queue_io_deq_bits_data;
  assign _T_783 = {{30'd0}, priority_0};
  assign _T_800 = _T_1931 & _T_754;
  assign _T_804 = _T_2228 & _T_758;
  assign _T_807 = _T_765[1:0];
  assign _T_808 = _T_812 == _T_807;
  assign _T_809 = _T_808 | reset;
  assign _T_811 = _T_809 == 1'h0;
  assign _T_812 = _T_765[1:0];
  assign _GEN_11 = 2'h1 == _T_807 ? enables_0_1 : enables_0_0;
  assign _GEN_12 = 2'h2 == _T_807 ? enables_0_2 : _GEN_11;
  assign _T_815 = _T_804 & _GEN_12;
  assign _T_832 = {{30'd0}, maxDevs_0};
  assign _T_853 = _T_2100 & _T_758;
  assign _GEN_13 = _T_853 ? _T_765 : {{30'd0}, priority_1};
  assign _T_872 = {{30'd0}, priority_1};
  assign _T_893 = _T_2108 & _T_758;
  assign _GEN_14 = _T_893 ? _T_765 : {{30'd0}, priority_2};
  assign _T_912 = {{30'd0}, priority_2};
  assign _T_933 = _T_2220 & _T_758;
  assign _GEN_15 = _T_933 ? _T_765 : {{30'd0}, threshold_0};
  assign _T_952 = {{30'd0}, threshold_0};
  assign _T_1013 = _T_2156 & _T_678;
  assign _GEN_17 = _T_1013 ? _T_685 : enables_0_1;
  assign _GEN_209 = {{1'd0}, enables_0_1};
  assign _T_1029 = _GEN_209 << 1;
  assign _GEN_210 = {{1'd0}, enables_0_0};
  assign _T_1033 = _GEN_210 | _T_1029;
  assign _T_1053 = _T_2156 & _T_718;
  assign _GEN_18 = _T_1053 ? _T_725 : enables_0_2;
  assign _GEN_211 = {{2'd0}, enables_0_2};
  assign _T_1069 = _GEN_211 << 2;
  assign _GEN_212 = {{1'd0}, _T_1033};
  assign _T_1073 = _GEN_212 | _T_1069;
  assign _T_1102 = Queue_io_deq_bits_index[0];
  assign _T_1103 = Queue_io_deq_bits_index[1];
  assign _T_1112 = Queue_io_deq_bits_index[10];
  assign _T_1113 = Queue_io_deq_bits_index[11];
  assign _T_1121 = Queue_io_deq_bits_index[19];
  assign _T_1126 = {_T_1103,_T_1102};
  assign _T_1127 = {_T_1121,_T_1113};
  assign _T_1128 = {_T_1127,_T_1112};
  assign _T_1129 = {_T_1128,_T_1126};
  assign _T_1165 = 32'h1 << _T_1129;
  assign _T_1167 = _T_1165[1];
  assign _T_1168 = _T_1165[2];
  assign _T_1174 = _T_1165[8];
  assign _T_1182 = _T_1165[16];
  assign _T_1183 = _T_1165[17];
  assign _T_1790 = Queue_io_deq_valid & io_tl_in_0_d_ready;
  assign _T_1791 = _T_1790 & Queue_io_deq_bits_read;
  assign _T_1930 = _T_1791 & _T_1183;
  assign _T_1931 = _T_1930 & _T_442;
  assign _T_2087 = Queue_io_deq_bits_read == 1'h0;
  assign _T_2088 = _T_1790 & _T_2087;
  assign _T_2099 = _T_2088 & _T_1167;
  assign _T_2100 = _T_2099 & _T_451;
  assign _T_2107 = _T_2088 & _T_1168;
  assign _T_2108 = _T_2107 & _T_460;
  assign _T_2155 = _T_2088 & _T_1174;
  assign _T_2156 = _T_2155 & _T_478;
  assign _T_2219 = _T_2088 & _T_1182;
  assign _T_2220 = _T_2219 & _T_469;
  assign _T_2227 = _T_2088 & _T_1183;
  assign _T_2228 = _T_2227 & _T_442;
  assign _T_2391 = Queue_io_deq_valid;
  assign _T_2432_4 = {{29'd0}, _T_744};
  assign _T_2432_8 = {{29'd0}, _T_1073};
  assign _GEN_143 = 5'h1 == _T_1129 ? _T_451 : _T_433;
  assign _GEN_144 = 5'h2 == _T_1129 ? _T_460 : _GEN_143;
  assign _GEN_145 = 5'h3 == _T_1129 ? 1'h1 : _GEN_144;
  assign _GEN_146 = 5'h4 == _T_1129 ? _T_424 : _GEN_145;
  assign _GEN_147 = 5'h5 == _T_1129 ? 1'h1 : _GEN_146;
  assign _GEN_148 = 5'h6 == _T_1129 ? 1'h1 : _GEN_147;
  assign _GEN_149 = 5'h7 == _T_1129 ? 1'h1 : _GEN_148;
  assign _GEN_150 = 5'h8 == _T_1129 ? _T_478 : _GEN_149;
  assign _GEN_151 = 5'h9 == _T_1129 ? 1'h1 : _GEN_150;
  assign _GEN_152 = 5'ha == _T_1129 ? 1'h1 : _GEN_151;
  assign _GEN_153 = 5'hb == _T_1129 ? 1'h1 : _GEN_152;
  assign _GEN_154 = 5'hc == _T_1129 ? 1'h1 : _GEN_153;
  assign _GEN_155 = 5'hd == _T_1129 ? 1'h1 : _GEN_154;
  assign _GEN_156 = 5'he == _T_1129 ? 1'h1 : _GEN_155;
  assign _GEN_157 = 5'hf == _T_1129 ? 1'h1 : _GEN_156;
  assign _GEN_158 = 5'h10 == _T_1129 ? _T_469 : _GEN_157;
  assign _GEN_159 = 5'h11 == _T_1129 ? _T_442 : _GEN_158;
  assign _GEN_160 = 5'h12 == _T_1129 ? 1'h1 : _GEN_159;
  assign _GEN_161 = 5'h13 == _T_1129 ? 1'h1 : _GEN_160;
  assign _GEN_162 = 5'h14 == _T_1129 ? 1'h1 : _GEN_161;
  assign _GEN_163 = 5'h15 == _T_1129 ? 1'h1 : _GEN_162;
  assign _GEN_164 = 5'h16 == _T_1129 ? 1'h1 : _GEN_163;
  assign _GEN_165 = 5'h17 == _T_1129 ? 1'h1 : _GEN_164;
  assign _GEN_166 = 5'h18 == _T_1129 ? 1'h1 : _GEN_165;
  assign _GEN_167 = 5'h19 == _T_1129 ? 1'h1 : _GEN_166;
  assign _GEN_168 = 5'h1a == _T_1129 ? 1'h1 : _GEN_167;
  assign _GEN_169 = 5'h1b == _T_1129 ? 1'h1 : _GEN_168;
  assign _GEN_170 = 5'h1c == _T_1129 ? 1'h1 : _GEN_169;
  assign _GEN_171 = 5'h1d == _T_1129 ? 1'h1 : _GEN_170;
  assign _GEN_172 = 5'h1e == _T_1129 ? 1'h1 : _GEN_171;
  assign _GEN_173 = 5'h1f == _T_1129 ? 1'h1 : _GEN_172;
  assign _GEN_174 = 5'h1 == _T_1129 ? _T_872 : _T_783;
  assign _GEN_175 = 5'h2 == _T_1129 ? _T_912 : _GEN_174;
  assign _GEN_176 = 5'h3 == _T_1129 ? 32'h0 : _GEN_175;
  assign _GEN_177 = 5'h4 == _T_1129 ? _T_2432_4 : _GEN_176;
  assign _GEN_178 = 5'h5 == _T_1129 ? 32'h0 : _GEN_177;
  assign _GEN_179 = 5'h6 == _T_1129 ? 32'h0 : _GEN_178;
  assign _GEN_180 = 5'h7 == _T_1129 ? 32'h0 : _GEN_179;
  assign _GEN_181 = 5'h8 == _T_1129 ? _T_2432_8 : _GEN_180;
  assign _GEN_182 = 5'h9 == _T_1129 ? 32'h0 : _GEN_181;
  assign _GEN_183 = 5'ha == _T_1129 ? 32'h0 : _GEN_182;
  assign _GEN_184 = 5'hb == _T_1129 ? 32'h0 : _GEN_183;
  assign _GEN_185 = 5'hc == _T_1129 ? 32'h0 : _GEN_184;
  assign _GEN_186 = 5'hd == _T_1129 ? 32'h0 : _GEN_185;
  assign _GEN_187 = 5'he == _T_1129 ? 32'h0 : _GEN_186;
  assign _GEN_188 = 5'hf == _T_1129 ? 32'h0 : _GEN_187;
  assign _GEN_189 = 5'h10 == _T_1129 ? _T_952 : _GEN_188;
  assign _GEN_190 = 5'h11 == _T_1129 ? _T_832 : _GEN_189;
  assign _GEN_191 = 5'h12 == _T_1129 ? 32'h0 : _GEN_190;
  assign _GEN_192 = 5'h13 == _T_1129 ? 32'h0 : _GEN_191;
  assign _GEN_193 = 5'h14 == _T_1129 ? 32'h0 : _GEN_192;
  assign _GEN_194 = 5'h15 == _T_1129 ? 32'h0 : _GEN_193;
  assign _GEN_195 = 5'h16 == _T_1129 ? 32'h0 : _GEN_194;
  assign _GEN_196 = 5'h17 == _T_1129 ? 32'h0 : _GEN_195;
  assign _GEN_197 = 5'h18 == _T_1129 ? 32'h0 : _GEN_196;
  assign _GEN_198 = 5'h19 == _T_1129 ? 32'h0 : _GEN_197;
  assign _GEN_199 = 5'h1a == _T_1129 ? 32'h0 : _GEN_198;
  assign _GEN_200 = 5'h1b == _T_1129 ? 32'h0 : _GEN_199;
  assign _GEN_201 = 5'h1c == _T_1129 ? 32'h0 : _GEN_200;
  assign _GEN_202 = 5'h1d == _T_1129 ? 32'h0 : _GEN_201;
  assign _GEN_203 = 5'h1e == _T_1129 ? 32'h0 : _GEN_202;
  assign _GEN_204 = 5'h1f == _T_1129 ? 32'h0 : _GEN_203;
  assign _T_2469 = _GEN_173 ? _GEN_204 : 32'h0;
  assign _T_2470 = _T_336_bits_extra[11:2];
  assign _T_2471 = _T_336_bits_extra[1:0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  priority_0 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  priority_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  priority_2 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  threshold_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  pending_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  pending_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  pending_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  enables_0_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  enables_0_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  enables_0_2 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  maxDevs_0 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_237 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    priority_0 <= 2'h0;
    priority_1 <= _GEN_13[1:0];
    priority_2 <= _GEN_14[1:0];
    threshold_0 <= _GEN_15[1:0];
    if (reset) begin
      pending_0 <= 1'h0;
    end else begin
      pending_0 <= 1'h0;
    end
    if (reset) begin
      pending_1 <= 1'h0;
    end else begin
      if (_T_285) begin
        pending_1 <= _T_287;
      end
    end
    if (reset) begin
      pending_2 <= 1'h0;
    end else begin
      if (_T_290) begin
        pending_2 <= _T_292;
      end
    end
    enables_0_0 <= 1'h0;
    if (_T_1013) begin
      enables_0_1 <= _T_685;
    end
    if (_T_1053) begin
      enables_0_2 <= _T_725;
    end
    if (_T_231) begin
      maxDevs_0 <= {{1'd0}, _T_229};
    end else begin
      maxDevs_0 <= 2'h2;
    end
    if (_T_231) begin
      if (_T_225) begin
        _T_237 <= 3'h4;
      end else begin
        _T_237 <= _T_220;
      end
    end else begin
      _T_237 <= _T_222;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_256) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Plic.scala:187 assert((claimer.asUInt & (claimer.asUInt - UInt(1))) === UInt(0)) // One-Hot\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_256) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_308) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Plic.scala:204 assert((completer.asUInt & (completer.asUInt - UInt(1))) === UInt(0)) // One-Hot\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_308) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_811) begin
          $fwrite(32'h80000002,"Assertion failed: completerDev should be consistent for all harts\n    at Plic.scala:220 assert(completerDev === data.extract(log2Ceil(nDevices+1)-1, 0),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_811) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CoreplexLocalInterrupter_clint(
  input         clock,
  input         reset,
  input         io_rtcTick,
  output        io_int_0_0,
  output        io_int_0_1,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [1:0]  io_in_0_a_bits_size,
  input  [9:0]  io_in_0_a_bits_source,
  input  [25:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [1:0]  io_in_0_d_bits_size,
  output [9:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error
);
  reg [31:0] time_0;
  reg [31:0] _RAND_0;
  reg [31:0] time_1;
  reg [31:0] _RAND_1;
  wire [63:0] _T_69;
  wire [64:0] _T_71;
  wire [63:0] _T_72;
  wire [31:0] _T_74;
  wire [63:0] _GEN_6;
  wire [31:0] _GEN_7;
  reg [31:0] timecmp_0_0;
  reg [31:0] _RAND_2;
  reg [31:0] timecmp_0_1;
  reg [31:0] _RAND_3;
  reg  ipi_0;
  reg [31:0] _RAND_4;
  wire [63:0] _T_81;
  wire  _T_82;
  wire [13:0] _T_88_bits_index;
  wire  _T_93;
  wire [23:0] _T_94;
  wire [11:0] _T_95;
  wire [13:0] _T_134;
  wire  _T_136;
  wire [13:0] _T_142;
  wire [13:0] _T_143;
  wire  _T_145;
  wire [13:0] _T_151;
  wire [13:0] _T_152;
  wire  _T_154;
  wire [13:0] _T_160;
  wire [13:0] _T_161;
  wire  _T_163;
  wire [13:0] _T_169;
  wire [13:0] _T_170;
  wire  _T_172;
  wire  _T_229;
  wire  _T_230;
  wire  _T_231;
  wire  _T_232;
  wire [7:0] _T_236;
  wire [7:0] _T_240;
  wire [7:0] _T_244;
  wire [7:0] _T_248;
  wire [15:0] _T_249;
  wire [15:0] _T_250;
  wire [31:0] _T_251;
  wire [31:0] _T_279;
  wire  _T_281;
  wire  _T_294;
  wire [31:0] _GEN_8;
  wire [31:0] _T_313;
  wire  _T_334;
  wire [31:0] _GEN_9;
  wire  _T_374;
  wire [63:0] _GEN_10;
  wire  _T_414;
  wire [31:0] _GEN_11;
  wire  _T_454;
  wire [31:0] _GEN_12;
  wire  _T_475;
  wire  _T_476;
  wire  _T_487;
  wire [1:0] _T_489;
  wire [2:0] _T_490;
  wire [7:0] _T_508;
  wire  _T_509;
  wire  _T_511;
  wire  _T_512;
  wire  _T_513;
  wire  _T_514;
  wire  _T_527;
  wire  _T_608;
  wire  _T_609;
  wire  _T_612;
  wire  _T_628;
  wire  _T_636;
  wire  _T_644;
  wire  _T_652;
  wire  _T_773;
  wire  _T_789;
  wire  _T_797;
  wire  _T_805;
  wire  _T_813;
  wire  _GEN_41;
  wire  _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire [31:0] _GEN_48;
  wire [31:0] _GEN_49;
  wire [31:0] _GEN_50;
  wire [31:0] _GEN_51;
  wire [31:0] _GEN_52;
  wire [31:0] _GEN_53;
  wire [31:0] _GEN_54;
  wire [31:0] _T_886;
  wire [9:0] _T_887;
  wire [1:0] _T_888;
  assign io_int_0_0 = ipi_0;
  assign io_int_0_1 = _T_82;
  assign io_in_0_a_ready = io_in_0_d_ready;
  assign io_in_0_d_valid = io_in_0_a_valid;
  assign io_in_0_d_bits_opcode = {{2'd0}, _T_93};
  assign io_in_0_d_bits_param = 2'h0;
  assign io_in_0_d_bits_size = _T_888;
  assign io_in_0_d_bits_source = _T_887;
  assign io_in_0_d_bits_sink = 1'h0;
  assign io_in_0_d_bits_data = _T_886;
  assign io_in_0_d_bits_error = 1'h0;
  assign _T_69 = {time_1,time_0};
  assign _T_71 = _T_69 + 64'h1;
  assign _T_72 = _T_71[63:0];
  assign _T_74 = _T_72[63:32];
  assign _GEN_6 = io_rtcTick ? _T_72 : {{32'd0}, time_0};
  assign _GEN_7 = io_rtcTick ? _T_74 : time_1;
  assign _T_81 = {timecmp_0_1,timecmp_0_0};
  assign _T_82 = _T_69 >= _T_81;
  assign _T_88_bits_index = _T_94[13:0];
  assign _T_93 = io_in_0_a_bits_opcode == 3'h4;
  assign _T_94 = io_in_0_a_bits_address[25:2];
  assign _T_95 = {io_in_0_a_bits_source,io_in_0_a_bits_size};
  assign _T_134 = _T_88_bits_index & 14'h2ffc;
  assign _T_136 = _T_134 == 14'h0;
  assign _T_142 = _T_88_bits_index ^ 14'h1001;
  assign _T_143 = _T_142 & 14'h2ffc;
  assign _T_145 = _T_143 == 14'h0;
  assign _T_151 = _T_88_bits_index ^ 14'h2ffe;
  assign _T_152 = _T_151 & 14'h2ffc;
  assign _T_154 = _T_152 == 14'h0;
  assign _T_160 = _T_88_bits_index ^ 14'h2fff;
  assign _T_161 = _T_160 & 14'h2ffc;
  assign _T_163 = _T_161 == 14'h0;
  assign _T_169 = _T_88_bits_index ^ 14'h1000;
  assign _T_170 = _T_169 & 14'h2ffc;
  assign _T_172 = _T_170 == 14'h0;
  assign _T_229 = io_in_0_a_bits_mask[0];
  assign _T_230 = io_in_0_a_bits_mask[1];
  assign _T_231 = io_in_0_a_bits_mask[2];
  assign _T_232 = io_in_0_a_bits_mask[3];
  assign _T_236 = _T_229 ? 8'hff : 8'h0;
  assign _T_240 = _T_230 ? 8'hff : 8'h0;
  assign _T_244 = _T_231 ? 8'hff : 8'h0;
  assign _T_248 = _T_232 ? 8'hff : 8'h0;
  assign _T_249 = {_T_240,_T_236};
  assign _T_250 = {_T_248,_T_244};
  assign _T_251 = {_T_250,_T_249};
  assign _T_279 = ~ _T_251;
  assign _T_281 = _T_279 == 32'h0;
  assign _T_294 = _T_773 & _T_281;
  assign _GEN_8 = _T_294 ? io_in_0_a_bits_data : {{31'd0}, ipi_0};
  assign _T_313 = {{31'd0}, ipi_0};
  assign _T_334 = _T_813 & _T_281;
  assign _GEN_9 = _T_334 ? io_in_0_a_bits_data : timecmp_0_1;
  assign _T_374 = _T_789 & _T_281;
  assign _GEN_10 = _T_374 ? {{32'd0}, io_in_0_a_bits_data} : _GEN_6;
  assign _T_414 = _T_797 & _T_281;
  assign _GEN_11 = _T_414 ? io_in_0_a_bits_data : _GEN_7;
  assign _T_454 = _T_805 & _T_281;
  assign _GEN_12 = _T_454 ? io_in_0_a_bits_data : timecmp_0_0;
  assign _T_475 = _T_88_bits_index[0];
  assign _T_476 = _T_88_bits_index[1];
  assign _T_487 = _T_88_bits_index[12];
  assign _T_489 = {_T_487,_T_476};
  assign _T_490 = {_T_489,_T_475};
  assign _T_508 = 8'h1 << _T_490;
  assign _T_509 = _T_508[0];
  assign _T_511 = _T_508[2];
  assign _T_512 = _T_508[3];
  assign _T_513 = _T_508[4];
  assign _T_514 = _T_508[5];
  assign _T_527 = io_in_0_a_valid & io_in_0_d_ready;
  assign _T_608 = _T_93 == 1'h0;
  assign _T_609 = _T_527 & _T_608;
  assign _T_612 = _T_609 & _T_509;
  assign _T_628 = _T_609 & _T_511;
  assign _T_636 = _T_609 & _T_512;
  assign _T_644 = _T_609 & _T_513;
  assign _T_652 = _T_609 & _T_514;
  assign _T_773 = _T_612 & _T_136;
  assign _T_789 = _T_628 & _T_154;
  assign _T_797 = _T_636 & _T_163;
  assign _T_805 = _T_644 & _T_172;
  assign _T_813 = _T_652 & _T_145;
  assign _GEN_41 = 3'h1 == _T_490 ? 1'h1 : _T_136;
  assign _GEN_42 = 3'h2 == _T_490 ? _T_154 : _GEN_41;
  assign _GEN_43 = 3'h3 == _T_490 ? _T_163 : _GEN_42;
  assign _GEN_44 = 3'h4 == _T_490 ? _T_172 : _GEN_43;
  assign _GEN_45 = 3'h5 == _T_490 ? _T_145 : _GEN_44;
  assign _GEN_46 = 3'h6 == _T_490 ? 1'h1 : _GEN_45;
  assign _GEN_47 = 3'h7 == _T_490 ? 1'h1 : _GEN_46;
  assign _GEN_48 = 3'h1 == _T_490 ? 32'h0 : _T_313;
  assign _GEN_49 = 3'h2 == _T_490 ? time_0 : _GEN_48;
  assign _GEN_50 = 3'h3 == _T_490 ? time_1 : _GEN_49;
  assign _GEN_51 = 3'h4 == _T_490 ? timecmp_0_0 : _GEN_50;
  assign _GEN_52 = 3'h5 == _T_490 ? timecmp_0_1 : _GEN_51;
  assign _GEN_53 = 3'h6 == _T_490 ? 32'h0 : _GEN_52;
  assign _GEN_54 = 3'h7 == _T_490 ? 32'h0 : _GEN_53;
  assign _T_886 = _GEN_47 ? _GEN_54 : 32'h0;
  assign _T_887 = _T_95[11:2];
  assign _T_888 = _T_95[1:0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  time_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  time_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  timecmp_0_0 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  timecmp_0_1 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  ipi_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      time_0 <= 32'h0;
    end else begin
      time_0 <= _GEN_10[31:0];
    end
    if (reset) begin
      time_1 <= 32'h0;
    end else begin
      if (_T_414) begin
        time_1 <= io_in_0_a_bits_data;
      end else begin
        if (io_rtcTick) begin
          time_1 <= _T_74;
        end
      end
    end
    if (_T_454) begin
      timecmp_0_0 <= io_in_0_a_bits_data;
    end
    if (_T_334) begin
      timecmp_0_1 <= io_in_0_a_bits_data;
    end
    if (reset) begin
      ipi_0 <= 1'h0;
    end else begin
      ipi_0 <= _GEN_8[0];
    end
  end
endmodule
module DMIToTL_dmi2tl(
  output        io_dmi_req_ready,
  input         io_dmi_req_valid,
  input  [6:0]  io_dmi_req_bits_addr,
  input  [31:0] io_dmi_req_bits_data,
  input  [1:0]  io_dmi_req_bits_op,
  input         io_dmi_resp_ready,
  output        io_dmi_resp_valid,
  output [31:0] io_dmi_resp_bits_data,
  output [1:0]  io_dmi_resp_bits_resp,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [1:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [8:0]  io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire [8:0] _GEN_21;
  wire [8:0] _T_57;
  wire  _T_203;
  wire  _T_205;
  wire  _T_207;
  wire  _T_208;
  wire [2:0] _GEN_7;
  wire [31:0] _GEN_13;
  wire  _T_212;
  wire  _T_213;
  wire [2:0] _GEN_14;
  wire [8:0] _GEN_18;
  wire [3:0] _GEN_19;
  wire [31:0] _GEN_20;
  assign io_dmi_req_ready = io_out_0_a_ready;
  assign io_dmi_resp_valid = io_out_0_d_valid;
  assign io_dmi_resp_bits_data = io_out_0_d_bits_data;
  assign io_dmi_resp_bits_resp = {{1'd0}, io_out_0_d_bits_error};
  assign io_out_0_a_valid = io_dmi_req_valid;
  assign io_out_0_a_bits_opcode = _GEN_14;
  assign io_out_0_a_bits_size = 2'h2;
  assign io_out_0_a_bits_source = 1'h0;
  assign io_out_0_a_bits_address = _GEN_18;
  assign io_out_0_a_bits_mask = _GEN_19;
  assign io_out_0_a_bits_data = _GEN_20;
  assign io_out_0_d_ready = io_dmi_resp_ready;
  assign _GEN_21 = {{2'd0}, io_dmi_req_bits_addr};
  assign _T_57 = _GEN_21 << 2;
  assign _T_203 = io_dmi_req_bits_op == 2'h2;
  assign _T_205 = io_dmi_req_bits_op == 2'h1;
  assign _T_207 = _T_203 == 1'h0;
  assign _T_208 = _T_207 & _T_205;
  assign _GEN_7 = _T_208 ? 3'h4 : 3'h0;
  assign _GEN_13 = _T_208 ? 32'h0 : io_dmi_req_bits_data;
  assign _T_212 = _T_205 == 1'h0;
  assign _T_213 = _T_207 & _T_212;
  assign _GEN_14 = _T_213 ? 3'h1 : _GEN_7;
  assign _GEN_18 = _T_213 ? 9'h40 : _T_57;
  assign _GEN_19 = _T_213 ? 4'h0 : 4'hf;
  assign _GEN_20 = _T_213 ? 32'h0 : _GEN_13;
endmodule
module TLXbar_dmiXbar(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [1:0]  io_in_0_a_bits_size,
  input         io_in_0_a_bits_source,
  input  [8:0]  io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_1_a_ready,
  output        io_out_1_a_valid,
  output [2:0]  io_out_1_a_bits_opcode,
  output [1:0]  io_out_1_a_bits_size,
  output        io_out_1_a_bits_source,
  output [8:0]  io_out_1_a_bits_address,
  output [3:0]  io_out_1_a_bits_mask,
  output [31:0] io_out_1_a_bits_data,
  output        io_out_1_d_ready,
  input         io_out_1_d_valid,
  input  [2:0]  io_out_1_d_bits_opcode,
  input  [1:0]  io_out_1_d_bits_param,
  input  [1:0]  io_out_1_d_bits_size,
  input         io_out_1_d_bits_source,
  input         io_out_1_d_bits_sink,
  input  [31:0] io_out_1_d_bits_data,
  input         io_out_1_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [1:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [6:0]  io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [1:0]  io_out_0_d_bits_size,
  input         io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire [8:0] _T_634;
  wire [9:0] _T_635;
  wire [9:0] _T_637;
  wire [9:0] _T_638;
  wire  _T_640;
  wire [9:0] _T_643;
  wire [9:0] _T_645;
  wire [9:0] _T_646;
  wire  _T_648;
  wire [8:0] _T_650;
  wire [9:0] _T_651;
  wire [9:0] _T_653;
  wire [9:0] _T_654;
  wire  _T_656;
  wire [8:0] _T_658;
  wire [9:0] _T_659;
  wire [9:0] _T_661;
  wire [9:0] _T_662;
  wire  _T_664;
  wire [8:0] _T_666;
  wire [9:0] _T_667;
  wire [9:0] _T_669;
  wire [9:0] _T_670;
  wire  _T_672;
  wire [8:0] _T_674;
  wire [9:0] _T_675;
  wire [9:0] _T_677;
  wire [9:0] _T_678;
  wire  _T_680;
  wire [8:0] _T_682;
  wire [9:0] _T_683;
  wire [9:0] _T_685;
  wire [9:0] _T_686;
  wire  _T_688;
  wire [8:0] _T_690;
  wire [9:0] _T_691;
  wire [9:0] _T_693;
  wire [9:0] _T_694;
  wire  _T_696;
  wire  _T_697;
  wire  _T_698;
  wire  _T_699;
  wire  _T_700;
  wire  _T_701;
  wire  _T_702;
  wire  _T_967;
  wire  _T_975;
  wire  _T_1226;
  wire  _T_1227;
  wire  _T_1230;
  wire  _T_1232;
  wire  _T_1233;
  wire  _T_1354;
  wire  _T_1379;
  wire  _T_1450;
  wire  _T_1457;
  wire  _T_1458;
  wire  _T_1460;
  wire  _T_1524;
  wire  _T_1531;
  wire  _T_1532;
  wire  _T_1534;
  reg  _T_1575;
  reg [31:0] _RAND_0;
  wire  _T_1577;
  wire  _T_1578;
  wire [1:0] _T_1579;
  wire  _T_1581;
  wire  _T_1582;
  wire  _T_1584;
  reg [1:0] _T_1588;
  reg [31:0] _RAND_1;
  wire [1:0] _T_1589;
  wire [1:0] _T_1590;
  wire [3:0] _T_1591;
  wire [2:0] _T_1592;
  wire [3:0] _GEN_1;
  wire [3:0] _T_1593;
  wire [2:0] _T_1595;
  wire [3:0] _GEN_2;
  wire [3:0] _T_1596;
  wire [3:0] _GEN_3;
  wire [3:0] _T_1597;
  wire [1:0] _T_1598;
  wire [1:0] _T_1599;
  wire [1:0] _T_1600;
  wire [1:0] _T_1601;
  wire  _T_1603;
  wire  _T_1604;
  wire [1:0] _T_1605;
  wire [2:0] _GEN_4;
  wire [2:0] _T_1606;
  wire [1:0] _T_1607;
  wire [1:0] _T_1608;
  wire [1:0] _GEN_0;
  wire  _T_1611;
  wire  _T_1612;
  wire  _T_1620;
  wire  _T_1621;
  wire  _T_1631;
  wire  _T_1635;
  wire  _T_1640;
  wire  _T_1641;
  wire  _T_1643;
  wire  _T_1645;
  wire  _T_1646;
  wire  _T_1648;
  wire  _T_1650;
  wire  _T_1651;
  wire  _T_1653;
  wire  _T_1659;
  wire [1:0] _T_1660;
  wire [1:0] _T_1661;
  wire  _T_1662;
  wire  _T_1663;
  reg  _T_1681_0;
  reg [31:0] _RAND_2;
  reg  _T_1681_1;
  reg [31:0] _RAND_3;
  wire  _T_1692_0;
  wire  _T_1692_1;
  wire  _T_1700_0;
  wire  _T_1700_1;
  wire  _T_1708;
  wire  _T_1709;
  wire  _T_1713;
  wire  _T_1715;
  wire  _T_1716;
  wire  _T_1719;
  wire [32:0] _T_1721;
  wire [33:0] _T_1722;
  wire [2:0] _T_1723;
  wire [4:0] _T_1724;
  wire [7:0] _T_1725;
  wire [41:0] _T_1726;
  wire [41:0] _T_1728;
  wire [32:0] _T_1729;
  wire [33:0] _T_1730;
  wire [2:0] _T_1731;
  wire [4:0] _T_1732;
  wire [7:0] _T_1733;
  wire [41:0] _T_1734;
  wire [41:0] _T_1736;
  wire [41:0] _T_1737;
  wire  _T_1742;
  wire [31:0] _T_1743;
  assign io_in_0_a_ready = _T_1233;
  assign io_in_0_d_valid = _T_1719;
  assign io_in_0_d_bits_data = _T_1743;
  assign io_in_0_d_bits_error = _T_1742;
  assign io_out_1_a_valid = _T_1227;
  assign io_out_1_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_1_a_bits_size = io_in_0_a_bits_size;
  assign io_out_1_a_bits_source = io_in_0_a_bits_source;
  assign io_out_1_a_bits_address = io_in_0_a_bits_address;
  assign io_out_1_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_1_a_bits_data = io_in_0_a_bits_data;
  assign io_out_1_d_ready = _T_1709;
  assign io_out_0_a_valid = _T_1226;
  assign io_out_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign io_out_0_a_bits_size = io_in_0_a_bits_size;
  assign io_out_0_a_bits_source = io_in_0_a_bits_source;
  assign io_out_0_a_bits_address = io_in_0_a_bits_address[6:0];
  assign io_out_0_a_bits_mask = io_in_0_a_bits_mask;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = _T_1708;
  assign _T_634 = io_in_0_a_bits_address ^ 9'h40;
  assign _T_635 = {1'b0,$signed(_T_634)};
  assign _T_637 = $signed(_T_635) & $signed(10'sh1fc);
  assign _T_638 = $signed(_T_637);
  assign _T_640 = $signed(_T_638) == $signed(10'sh0);
  assign _T_643 = {1'b0,$signed(io_in_0_a_bits_address)};
  assign _T_645 = $signed(_T_643) & $signed(10'sh1c0);
  assign _T_646 = $signed(_T_645);
  assign _T_648 = $signed(_T_646) == $signed(10'sh0);
  assign _T_650 = io_in_0_a_bits_address ^ 9'h44;
  assign _T_651 = {1'b0,$signed(_T_650)};
  assign _T_653 = $signed(_T_651) & $signed(10'sh1fc);
  assign _T_654 = $signed(_T_653);
  assign _T_656 = $signed(_T_654) == $signed(10'sh0);
  assign _T_658 = io_in_0_a_bits_address ^ 9'h48;
  assign _T_659 = {1'b0,$signed(_T_658)};
  assign _T_661 = $signed(_T_659) & $signed(10'sh1f8);
  assign _T_662 = $signed(_T_661);
  assign _T_664 = $signed(_T_662) == $signed(10'sh0);
  assign _T_666 = io_in_0_a_bits_address ^ 9'h50;
  assign _T_667 = {1'b0,$signed(_T_666)};
  assign _T_669 = $signed(_T_667) & $signed(10'sh1f0);
  assign _T_670 = $signed(_T_669);
  assign _T_672 = $signed(_T_670) == $signed(10'sh0);
  assign _T_674 = io_in_0_a_bits_address ^ 9'h60;
  assign _T_675 = {1'b0,$signed(_T_674)};
  assign _T_677 = $signed(_T_675) & $signed(10'sh1e0);
  assign _T_678 = $signed(_T_677);
  assign _T_680 = $signed(_T_678) == $signed(10'sh0);
  assign _T_682 = io_in_0_a_bits_address ^ 9'h80;
  assign _T_683 = {1'b0,$signed(_T_682)};
  assign _T_685 = $signed(_T_683) & $signed(10'sh180);
  assign _T_686 = $signed(_T_685);
  assign _T_688 = $signed(_T_686) == $signed(10'sh0);
  assign _T_690 = io_in_0_a_bits_address ^ 9'h100;
  assign _T_691 = {1'b0,$signed(_T_690)};
  assign _T_693 = $signed(_T_691) & $signed(10'sh100);
  assign _T_694 = $signed(_T_693);
  assign _T_696 = $signed(_T_694) == $signed(10'sh0);
  assign _T_697 = _T_648 | _T_656;
  assign _T_698 = _T_697 | _T_664;
  assign _T_699 = _T_698 | _T_672;
  assign _T_700 = _T_699 | _T_680;
  assign _T_701 = _T_700 | _T_688;
  assign _T_702 = _T_701 | _T_696;
  assign _T_967 = io_out_0_d_bits_source == 1'h0;
  assign _T_975 = io_out_1_d_bits_source == 1'h0;
  assign _T_1226 = io_in_0_a_valid & _T_640;
  assign _T_1227 = io_in_0_a_valid & _T_702;
  assign _T_1230 = _T_640 ? io_out_0_a_ready : 1'h0;
  assign _T_1232 = _T_702 ? io_out_1_a_ready : 1'h0;
  assign _T_1233 = _T_1230 | _T_1232;
  assign _T_1354 = io_out_0_d_valid & _T_967;
  assign _T_1379 = io_out_1_d_valid & _T_975;
  assign _T_1450 = _T_1226 == 1'h0;
  assign _T_1457 = _T_1450 | _T_1226;
  assign _T_1458 = _T_1457 | reset;
  assign _T_1460 = _T_1458 == 1'h0;
  assign _T_1524 = _T_1227 == 1'h0;
  assign _T_1531 = _T_1524 | _T_1227;
  assign _T_1532 = _T_1531 | reset;
  assign _T_1534 = _T_1532 == 1'h0;
  assign _T_1577 = _T_1575 == 1'h0;
  assign _T_1578 = _T_1577 & io_in_0_d_ready;
  assign _T_1579 = {_T_1379,_T_1354};
  assign _T_1581 = _T_1579 == _T_1579;
  assign _T_1582 = _T_1581 | reset;
  assign _T_1584 = _T_1582 == 1'h0;
  assign _T_1589 = ~ _T_1588;
  assign _T_1590 = _T_1579 & _T_1589;
  assign _T_1591 = {_T_1590,_T_1579};
  assign _T_1592 = _T_1591[3:1];
  assign _GEN_1 = {{1'd0}, _T_1592};
  assign _T_1593 = _T_1591 | _GEN_1;
  assign _T_1595 = _T_1593[3:1];
  assign _GEN_2 = {{2'd0}, _T_1588};
  assign _T_1596 = _GEN_2 << 2;
  assign _GEN_3 = {{1'd0}, _T_1595};
  assign _T_1597 = _GEN_3 | _T_1596;
  assign _T_1598 = _T_1597[3:2];
  assign _T_1599 = _T_1597[1:0];
  assign _T_1600 = _T_1598 & _T_1599;
  assign _T_1601 = ~ _T_1600;
  assign _T_1603 = _T_1579 != 2'h0;
  assign _T_1604 = _T_1578 & _T_1603;
  assign _T_1605 = _T_1601 & _T_1579;
  assign _GEN_4 = {{1'd0}, _T_1605};
  assign _T_1606 = _GEN_4 << 1;
  assign _T_1607 = _T_1606[1:0];
  assign _T_1608 = _T_1605 | _T_1607;
  assign _GEN_0 = _T_1604 ? _T_1608 : _T_1588;
  assign _T_1611 = _T_1601[0];
  assign _T_1612 = _T_1601[1];
  assign _T_1620 = _T_1611 & _T_1354;
  assign _T_1621 = _T_1612 & _T_1379;
  assign _T_1631 = _T_1620 | _T_1621;
  assign _T_1635 = _T_1620 == 1'h0;
  assign _T_1640 = _T_1621 == 1'h0;
  assign _T_1641 = _T_1635 | _T_1640;
  assign _T_1643 = _T_1641 | reset;
  assign _T_1645 = _T_1643 == 1'h0;
  assign _T_1646 = _T_1354 | _T_1379;
  assign _T_1648 = _T_1646 == 1'h0;
  assign _T_1650 = _T_1648 | _T_1631;
  assign _T_1651 = _T_1650 | reset;
  assign _T_1653 = _T_1651 == 1'h0;
  assign _T_1659 = io_in_0_d_ready & _T_1719;
  assign _T_1660 = _T_1575 - _T_1659;
  assign _T_1661 = $unsigned(_T_1660);
  assign _T_1662 = _T_1661[0:0];
  assign _T_1663 = _T_1578 ? 1'h0 : _T_1662;
  assign _T_1692_0 = _T_1577 ? _T_1620 : _T_1681_0;
  assign _T_1692_1 = _T_1577 ? _T_1621 : _T_1681_1;
  assign _T_1700_0 = _T_1577 ? _T_1611 : _T_1681_0;
  assign _T_1700_1 = _T_1577 ? _T_1612 : _T_1681_1;
  assign _T_1708 = io_in_0_d_ready & _T_1700_0;
  assign _T_1709 = io_in_0_d_ready & _T_1700_1;
  assign _T_1713 = _T_1681_0 ? _T_1354 : 1'h0;
  assign _T_1715 = _T_1681_1 ? _T_1379 : 1'h0;
  assign _T_1716 = _T_1713 | _T_1715;
  assign _T_1719 = _T_1577 ? _T_1646 : _T_1716;
  assign _T_1721 = {io_out_0_d_bits_sink,io_out_0_d_bits_data};
  assign _T_1722 = {_T_1721,io_out_0_d_bits_error};
  assign _T_1723 = {io_out_0_d_bits_size,io_out_0_d_bits_source};
  assign _T_1724 = {io_out_0_d_bits_opcode,io_out_0_d_bits_param};
  assign _T_1725 = {_T_1724,_T_1723};
  assign _T_1726 = {_T_1725,_T_1722};
  assign _T_1728 = _T_1692_0 ? _T_1726 : 42'h0;
  assign _T_1729 = {io_out_1_d_bits_sink,io_out_1_d_bits_data};
  assign _T_1730 = {_T_1729,io_out_1_d_bits_error};
  assign _T_1731 = {io_out_1_d_bits_size,io_out_1_d_bits_source};
  assign _T_1732 = {io_out_1_d_bits_opcode,io_out_1_d_bits_param};
  assign _T_1733 = {_T_1732,_T_1731};
  assign _T_1734 = {_T_1733,_T_1730};
  assign _T_1736 = _T_1692_1 ? _T_1734 : 42'h0;
  assign _T_1737 = _T_1728 | _T_1736;
  assign _T_1742 = _T_1737[0];
  assign _T_1743 = _T_1737[32:1];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1575 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1588 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_1681_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_1681_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1575 <= 1'h0;
    end else begin
      if (_T_1578) begin
        _T_1575 <= 1'h0;
      end else begin
        _T_1575 <= _T_1662;
      end
    end
    if (reset) begin
      _T_1588 <= 2'h3;
    end else begin
      if (_T_1604) begin
        _T_1588 <= _T_1608;
      end
    end
    if (reset) begin
      _T_1681_0 <= 1'h0;
    end else begin
      if (_T_1577) begin
        _T_1681_0 <= _T_1620;
      end
    end
    if (reset) begin
      _T_1681_1 <= 1'h0;
    end else begin
      if (_T_1577) begin
        _T_1681_1 <= _T_1621;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1460) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1460) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1534) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1534) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1584) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1584) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1645) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1645) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AsyncResetRegVec(
  input         clock,
  input         reset,
  input  [31:0] io_d,
  output [31:0] io_q,
  input         io_en
);
  wire  reg_0_rst;
  wire  reg_0_clk;
  wire  reg_0_en;
  wire  reg_0_q;
  wire  reg_0_d;
  wire  reg_1_rst;
  wire  reg_1_clk;
  wire  reg_1_en;
  wire  reg_1_q;
  wire  reg_1_d;
  wire  reg_2_rst;
  wire  reg_2_clk;
  wire  reg_2_en;
  wire  reg_2_q;
  wire  reg_2_d;
  wire  reg_3_rst;
  wire  reg_3_clk;
  wire  reg_3_en;
  wire  reg_3_q;
  wire  reg_3_d;
  wire  reg_4_rst;
  wire  reg_4_clk;
  wire  reg_4_en;
  wire  reg_4_q;
  wire  reg_4_d;
  wire  reg_5_rst;
  wire  reg_5_clk;
  wire  reg_5_en;
  wire  reg_5_q;
  wire  reg_5_d;
  wire  reg_6_rst;
  wire  reg_6_clk;
  wire  reg_6_en;
  wire  reg_6_q;
  wire  reg_6_d;
  wire  reg_7_rst;
  wire  reg_7_clk;
  wire  reg_7_en;
  wire  reg_7_q;
  wire  reg_7_d;
  wire  reg_8_rst;
  wire  reg_8_clk;
  wire  reg_8_en;
  wire  reg_8_q;
  wire  reg_8_d;
  wire  reg_9_rst;
  wire  reg_9_clk;
  wire  reg_9_en;
  wire  reg_9_q;
  wire  reg_9_d;
  wire  reg_10_rst;
  wire  reg_10_clk;
  wire  reg_10_en;
  wire  reg_10_q;
  wire  reg_10_d;
  wire  reg_11_rst;
  wire  reg_11_clk;
  wire  reg_11_en;
  wire  reg_11_q;
  wire  reg_11_d;
  wire  reg_12_rst;
  wire  reg_12_clk;
  wire  reg_12_en;
  wire  reg_12_q;
  wire  reg_12_d;
  wire  reg_13_rst;
  wire  reg_13_clk;
  wire  reg_13_en;
  wire  reg_13_q;
  wire  reg_13_d;
  wire  reg_14_rst;
  wire  reg_14_clk;
  wire  reg_14_en;
  wire  reg_14_q;
  wire  reg_14_d;
  wire  reg_15_rst;
  wire  reg_15_clk;
  wire  reg_15_en;
  wire  reg_15_q;
  wire  reg_15_d;
  wire  reg_16_rst;
  wire  reg_16_clk;
  wire  reg_16_en;
  wire  reg_16_q;
  wire  reg_16_d;
  wire  reg_17_rst;
  wire  reg_17_clk;
  wire  reg_17_en;
  wire  reg_17_q;
  wire  reg_17_d;
  wire  reg_18_rst;
  wire  reg_18_clk;
  wire  reg_18_en;
  wire  reg_18_q;
  wire  reg_18_d;
  wire  reg_19_rst;
  wire  reg_19_clk;
  wire  reg_19_en;
  wire  reg_19_q;
  wire  reg_19_d;
  wire  reg_20_rst;
  wire  reg_20_clk;
  wire  reg_20_en;
  wire  reg_20_q;
  wire  reg_20_d;
  wire  reg_21_rst;
  wire  reg_21_clk;
  wire  reg_21_en;
  wire  reg_21_q;
  wire  reg_21_d;
  wire  reg_22_rst;
  wire  reg_22_clk;
  wire  reg_22_en;
  wire  reg_22_q;
  wire  reg_22_d;
  wire  reg_23_rst;
  wire  reg_23_clk;
  wire  reg_23_en;
  wire  reg_23_q;
  wire  reg_23_d;
  wire  reg_24_rst;
  wire  reg_24_clk;
  wire  reg_24_en;
  wire  reg_24_q;
  wire  reg_24_d;
  wire  reg_25_rst;
  wire  reg_25_clk;
  wire  reg_25_en;
  wire  reg_25_q;
  wire  reg_25_d;
  wire  reg_26_rst;
  wire  reg_26_clk;
  wire  reg_26_en;
  wire  reg_26_q;
  wire  reg_26_d;
  wire  reg_27_rst;
  wire  reg_27_clk;
  wire  reg_27_en;
  wire  reg_27_q;
  wire  reg_27_d;
  wire  reg_28_rst;
  wire  reg_28_clk;
  wire  reg_28_en;
  wire  reg_28_q;
  wire  reg_28_d;
  wire  reg_29_rst;
  wire  reg_29_clk;
  wire  reg_29_en;
  wire  reg_29_q;
  wire  reg_29_d;
  wire  reg_30_rst;
  wire  reg_30_clk;
  wire  reg_30_en;
  wire  reg_30_q;
  wire  reg_30_d;
  wire  reg_31_rst;
  wire  reg_31_clk;
  wire  reg_31_en;
  wire  reg_31_q;
  wire  reg_31_d;
  wire  _T_5;
  wire  _T_6;
  wire  _T_7;
  wire  _T_8;
  wire  _T_9;
  wire  _T_10;
  wire  _T_11;
  wire  _T_12;
  wire  _T_13;
  wire  _T_14;
  wire  _T_15;
  wire  _T_16;
  wire  _T_17;
  wire  _T_18;
  wire  _T_19;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_36;
  wire [1:0] _T_37;
  wire [1:0] _T_38;
  wire [3:0] _T_39;
  wire [1:0] _T_40;
  wire [1:0] _T_41;
  wire [3:0] _T_42;
  wire [7:0] _T_43;
  wire [1:0] _T_44;
  wire [1:0] _T_45;
  wire [3:0] _T_46;
  wire [1:0] _T_47;
  wire [1:0] _T_48;
  wire [3:0] _T_49;
  wire [7:0] _T_50;
  wire [15:0] _T_51;
  wire [1:0] _T_52;
  wire [1:0] _T_53;
  wire [3:0] _T_54;
  wire [1:0] _T_55;
  wire [1:0] _T_56;
  wire [3:0] _T_57;
  wire [7:0] _T_58;
  wire [1:0] _T_59;
  wire [1:0] _T_60;
  wire [3:0] _T_61;
  wire [1:0] _T_62;
  wire [1:0] _T_63;
  wire [3:0] _T_64;
  wire [7:0] _T_65;
  wire [15:0] _T_66;
  wire [31:0] _T_67;
  AsyncResetReg reg_0 (
    .rst(reg_0_rst),
    .clk(reg_0_clk),
    .en(reg_0_en),
    .q(reg_0_q),
    .d(reg_0_d)
  );
  AsyncResetReg reg_1 (
    .rst(reg_1_rst),
    .clk(reg_1_clk),
    .en(reg_1_en),
    .q(reg_1_q),
    .d(reg_1_d)
  );
  AsyncResetReg reg_2 (
    .rst(reg_2_rst),
    .clk(reg_2_clk),
    .en(reg_2_en),
    .q(reg_2_q),
    .d(reg_2_d)
  );
  AsyncResetReg reg_3 (
    .rst(reg_3_rst),
    .clk(reg_3_clk),
    .en(reg_3_en),
    .q(reg_3_q),
    .d(reg_3_d)
  );
  AsyncResetReg reg_4 (
    .rst(reg_4_rst),
    .clk(reg_4_clk),
    .en(reg_4_en),
    .q(reg_4_q),
    .d(reg_4_d)
  );
  AsyncResetReg reg_5 (
    .rst(reg_5_rst),
    .clk(reg_5_clk),
    .en(reg_5_en),
    .q(reg_5_q),
    .d(reg_5_d)
  );
  AsyncResetReg reg_6 (
    .rst(reg_6_rst),
    .clk(reg_6_clk),
    .en(reg_6_en),
    .q(reg_6_q),
    .d(reg_6_d)
  );
  AsyncResetReg reg_7 (
    .rst(reg_7_rst),
    .clk(reg_7_clk),
    .en(reg_7_en),
    .q(reg_7_q),
    .d(reg_7_d)
  );
  AsyncResetReg reg_8 (
    .rst(reg_8_rst),
    .clk(reg_8_clk),
    .en(reg_8_en),
    .q(reg_8_q),
    .d(reg_8_d)
  );
  AsyncResetReg reg_9 (
    .rst(reg_9_rst),
    .clk(reg_9_clk),
    .en(reg_9_en),
    .q(reg_9_q),
    .d(reg_9_d)
  );
  AsyncResetReg reg_10 (
    .rst(reg_10_rst),
    .clk(reg_10_clk),
    .en(reg_10_en),
    .q(reg_10_q),
    .d(reg_10_d)
  );
  AsyncResetReg reg_11 (
    .rst(reg_11_rst),
    .clk(reg_11_clk),
    .en(reg_11_en),
    .q(reg_11_q),
    .d(reg_11_d)
  );
  AsyncResetReg reg_12 (
    .rst(reg_12_rst),
    .clk(reg_12_clk),
    .en(reg_12_en),
    .q(reg_12_q),
    .d(reg_12_d)
  );
  AsyncResetReg reg_13 (
    .rst(reg_13_rst),
    .clk(reg_13_clk),
    .en(reg_13_en),
    .q(reg_13_q),
    .d(reg_13_d)
  );
  AsyncResetReg reg_14 (
    .rst(reg_14_rst),
    .clk(reg_14_clk),
    .en(reg_14_en),
    .q(reg_14_q),
    .d(reg_14_d)
  );
  AsyncResetReg reg_15 (
    .rst(reg_15_rst),
    .clk(reg_15_clk),
    .en(reg_15_en),
    .q(reg_15_q),
    .d(reg_15_d)
  );
  AsyncResetReg reg_16 (
    .rst(reg_16_rst),
    .clk(reg_16_clk),
    .en(reg_16_en),
    .q(reg_16_q),
    .d(reg_16_d)
  );
  AsyncResetReg reg_17 (
    .rst(reg_17_rst),
    .clk(reg_17_clk),
    .en(reg_17_en),
    .q(reg_17_q),
    .d(reg_17_d)
  );
  AsyncResetReg reg_18 (
    .rst(reg_18_rst),
    .clk(reg_18_clk),
    .en(reg_18_en),
    .q(reg_18_q),
    .d(reg_18_d)
  );
  AsyncResetReg reg_19 (
    .rst(reg_19_rst),
    .clk(reg_19_clk),
    .en(reg_19_en),
    .q(reg_19_q),
    .d(reg_19_d)
  );
  AsyncResetReg reg_20 (
    .rst(reg_20_rst),
    .clk(reg_20_clk),
    .en(reg_20_en),
    .q(reg_20_q),
    .d(reg_20_d)
  );
  AsyncResetReg reg_21 (
    .rst(reg_21_rst),
    .clk(reg_21_clk),
    .en(reg_21_en),
    .q(reg_21_q),
    .d(reg_21_d)
  );
  AsyncResetReg reg_22 (
    .rst(reg_22_rst),
    .clk(reg_22_clk),
    .en(reg_22_en),
    .q(reg_22_q),
    .d(reg_22_d)
  );
  AsyncResetReg reg_23 (
    .rst(reg_23_rst),
    .clk(reg_23_clk),
    .en(reg_23_en),
    .q(reg_23_q),
    .d(reg_23_d)
  );
  AsyncResetReg reg_24 (
    .rst(reg_24_rst),
    .clk(reg_24_clk),
    .en(reg_24_en),
    .q(reg_24_q),
    .d(reg_24_d)
  );
  AsyncResetReg reg_25 (
    .rst(reg_25_rst),
    .clk(reg_25_clk),
    .en(reg_25_en),
    .q(reg_25_q),
    .d(reg_25_d)
  );
  AsyncResetReg reg_26 (
    .rst(reg_26_rst),
    .clk(reg_26_clk),
    .en(reg_26_en),
    .q(reg_26_q),
    .d(reg_26_d)
  );
  AsyncResetReg reg_27 (
    .rst(reg_27_rst),
    .clk(reg_27_clk),
    .en(reg_27_en),
    .q(reg_27_q),
    .d(reg_27_d)
  );
  AsyncResetReg reg_28 (
    .rst(reg_28_rst),
    .clk(reg_28_clk),
    .en(reg_28_en),
    .q(reg_28_q),
    .d(reg_28_d)
  );
  AsyncResetReg reg_29 (
    .rst(reg_29_rst),
    .clk(reg_29_clk),
    .en(reg_29_en),
    .q(reg_29_q),
    .d(reg_29_d)
  );
  AsyncResetReg reg_30 (
    .rst(reg_30_rst),
    .clk(reg_30_clk),
    .en(reg_30_en),
    .q(reg_30_q),
    .d(reg_30_d)
  );
  AsyncResetReg reg_31 (
    .rst(reg_31_rst),
    .clk(reg_31_clk),
    .en(reg_31_en),
    .q(reg_31_q),
    .d(reg_31_d)
  );
  assign io_q = _T_67;
  assign reg_0_rst = reset;
  assign reg_0_clk = clock;
  assign reg_0_en = io_en;
  assign reg_0_d = _T_5;
  assign reg_1_rst = reset;
  assign reg_1_clk = clock;
  assign reg_1_en = io_en;
  assign reg_1_d = _T_6;
  assign reg_2_rst = reset;
  assign reg_2_clk = clock;
  assign reg_2_en = io_en;
  assign reg_2_d = _T_7;
  assign reg_3_rst = reset;
  assign reg_3_clk = clock;
  assign reg_3_en = io_en;
  assign reg_3_d = _T_8;
  assign reg_4_rst = reset;
  assign reg_4_clk = clock;
  assign reg_4_en = io_en;
  assign reg_4_d = _T_9;
  assign reg_5_rst = reset;
  assign reg_5_clk = clock;
  assign reg_5_en = io_en;
  assign reg_5_d = _T_10;
  assign reg_6_rst = reset;
  assign reg_6_clk = clock;
  assign reg_6_en = io_en;
  assign reg_6_d = _T_11;
  assign reg_7_rst = reset;
  assign reg_7_clk = clock;
  assign reg_7_en = io_en;
  assign reg_7_d = _T_12;
  assign reg_8_rst = reset;
  assign reg_8_clk = clock;
  assign reg_8_en = io_en;
  assign reg_8_d = _T_13;
  assign reg_9_rst = reset;
  assign reg_9_clk = clock;
  assign reg_9_en = io_en;
  assign reg_9_d = _T_14;
  assign reg_10_rst = reset;
  assign reg_10_clk = clock;
  assign reg_10_en = io_en;
  assign reg_10_d = _T_15;
  assign reg_11_rst = reset;
  assign reg_11_clk = clock;
  assign reg_11_en = io_en;
  assign reg_11_d = _T_16;
  assign reg_12_rst = reset;
  assign reg_12_clk = clock;
  assign reg_12_en = io_en;
  assign reg_12_d = _T_17;
  assign reg_13_rst = reset;
  assign reg_13_clk = clock;
  assign reg_13_en = io_en;
  assign reg_13_d = _T_18;
  assign reg_14_rst = reset;
  assign reg_14_clk = clock;
  assign reg_14_en = io_en;
  assign reg_14_d = _T_19;
  assign reg_15_rst = reset;
  assign reg_15_clk = clock;
  assign reg_15_en = io_en;
  assign reg_15_d = _T_20;
  assign reg_16_rst = reset;
  assign reg_16_clk = clock;
  assign reg_16_en = io_en;
  assign reg_16_d = _T_21;
  assign reg_17_rst = reset;
  assign reg_17_clk = clock;
  assign reg_17_en = io_en;
  assign reg_17_d = _T_22;
  assign reg_18_rst = reset;
  assign reg_18_clk = clock;
  assign reg_18_en = io_en;
  assign reg_18_d = _T_23;
  assign reg_19_rst = reset;
  assign reg_19_clk = clock;
  assign reg_19_en = io_en;
  assign reg_19_d = _T_24;
  assign reg_20_rst = reset;
  assign reg_20_clk = clock;
  assign reg_20_en = io_en;
  assign reg_20_d = _T_25;
  assign reg_21_rst = reset;
  assign reg_21_clk = clock;
  assign reg_21_en = io_en;
  assign reg_21_d = _T_26;
  assign reg_22_rst = reset;
  assign reg_22_clk = clock;
  assign reg_22_en = io_en;
  assign reg_22_d = _T_27;
  assign reg_23_rst = reset;
  assign reg_23_clk = clock;
  assign reg_23_en = io_en;
  assign reg_23_d = _T_28;
  assign reg_24_rst = reset;
  assign reg_24_clk = clock;
  assign reg_24_en = io_en;
  assign reg_24_d = _T_29;
  assign reg_25_rst = reset;
  assign reg_25_clk = clock;
  assign reg_25_en = io_en;
  assign reg_25_d = _T_30;
  assign reg_26_rst = reset;
  assign reg_26_clk = clock;
  assign reg_26_en = io_en;
  assign reg_26_d = _T_31;
  assign reg_27_rst = reset;
  assign reg_27_clk = clock;
  assign reg_27_en = io_en;
  assign reg_27_d = _T_32;
  assign reg_28_rst = reset;
  assign reg_28_clk = clock;
  assign reg_28_en = io_en;
  assign reg_28_d = _T_33;
  assign reg_29_rst = reset;
  assign reg_29_clk = clock;
  assign reg_29_en = io_en;
  assign reg_29_d = _T_34;
  assign reg_30_rst = reset;
  assign reg_30_clk = clock;
  assign reg_30_en = io_en;
  assign reg_30_d = _T_35;
  assign reg_31_rst = reset;
  assign reg_31_clk = clock;
  assign reg_31_en = io_en;
  assign reg_31_d = _T_36;
  assign _T_5 = io_d[0];
  assign _T_6 = io_d[1];
  assign _T_7 = io_d[2];
  assign _T_8 = io_d[3];
  assign _T_9 = io_d[4];
  assign _T_10 = io_d[5];
  assign _T_11 = io_d[6];
  assign _T_12 = io_d[7];
  assign _T_13 = io_d[8];
  assign _T_14 = io_d[9];
  assign _T_15 = io_d[10];
  assign _T_16 = io_d[11];
  assign _T_17 = io_d[12];
  assign _T_18 = io_d[13];
  assign _T_19 = io_d[14];
  assign _T_20 = io_d[15];
  assign _T_21 = io_d[16];
  assign _T_22 = io_d[17];
  assign _T_23 = io_d[18];
  assign _T_24 = io_d[19];
  assign _T_25 = io_d[20];
  assign _T_26 = io_d[21];
  assign _T_27 = io_d[22];
  assign _T_28 = io_d[23];
  assign _T_29 = io_d[24];
  assign _T_30 = io_d[25];
  assign _T_31 = io_d[26];
  assign _T_32 = io_d[27];
  assign _T_33 = io_d[28];
  assign _T_34 = io_d[29];
  assign _T_35 = io_d[30];
  assign _T_36 = io_d[31];
  assign _T_37 = {reg_1_q,reg_0_q};
  assign _T_38 = {reg_3_q,reg_2_q};
  assign _T_39 = {_T_38,_T_37};
  assign _T_40 = {reg_5_q,reg_4_q};
  assign _T_41 = {reg_7_q,reg_6_q};
  assign _T_42 = {_T_41,_T_40};
  assign _T_43 = {_T_42,_T_39};
  assign _T_44 = {reg_9_q,reg_8_q};
  assign _T_45 = {reg_11_q,reg_10_q};
  assign _T_46 = {_T_45,_T_44};
  assign _T_47 = {reg_13_q,reg_12_q};
  assign _T_48 = {reg_15_q,reg_14_q};
  assign _T_49 = {_T_48,_T_47};
  assign _T_50 = {_T_49,_T_46};
  assign _T_51 = {_T_50,_T_43};
  assign _T_52 = {reg_17_q,reg_16_q};
  assign _T_53 = {reg_19_q,reg_18_q};
  assign _T_54 = {_T_53,_T_52};
  assign _T_55 = {reg_21_q,reg_20_q};
  assign _T_56 = {reg_23_q,reg_22_q};
  assign _T_57 = {_T_56,_T_55};
  assign _T_58 = {_T_57,_T_54};
  assign _T_59 = {reg_25_q,reg_24_q};
  assign _T_60 = {reg_27_q,reg_26_q};
  assign _T_61 = {_T_60,_T_59};
  assign _T_62 = {reg_29_q,reg_28_q};
  assign _T_63 = {reg_31_q,reg_30_q};
  assign _T_64 = {_T_63,_T_62};
  assign _T_65 = {_T_64,_T_61};
  assign _T_66 = {_T_65,_T_58};
  assign _T_67 = {_T_66,_T_51};
endmodule
module AsyncResetRegVec_1(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q,
  input   io_en
);
  wire  reg_0_rst;
  wire  reg_0_clk;
  wire  reg_0_en;
  wire  reg_0_q;
  wire  reg_0_d;
  AsyncResetReg reg_0 (
    .rst(reg_0_rst),
    .clk(reg_0_clk),
    .en(reg_0_en),
    .q(reg_0_q),
    .d(reg_0_d)
  );
  assign io_q = reg_0_q;
  assign reg_0_rst = reset;
  assign reg_0_clk = clock;
  assign reg_0_en = io_en;
  assign reg_0_d = io_d;
endmodule
module TLDebugModuleOuter_dmOuter(
  input         clock,
  input         reset,
  output        io_debugInterrupts_0_0,
  output        io_ctrl_ndreset,
  output        io_ctrl_dmactive,
  output        io_tlIn_0_a_ready,
  input         io_tlIn_0_a_valid,
  input  [2:0]  io_tlIn_0_a_bits_opcode,
  input  [1:0]  io_tlIn_0_a_bits_size,
  input         io_tlIn_0_a_bits_source,
  input  [6:0]  io_tlIn_0_a_bits_address,
  input  [3:0]  io_tlIn_0_a_bits_mask,
  input  [31:0] io_tlIn_0_a_bits_data,
  input         io_tlIn_0_d_ready,
  output        io_tlIn_0_d_valid,
  output [2:0]  io_tlIn_0_d_bits_opcode,
  output [1:0]  io_tlIn_0_d_bits_param,
  output [1:0]  io_tlIn_0_d_bits_size,
  output        io_tlIn_0_d_bits_source,
  output        io_tlIn_0_d_bits_sink,
  output [31:0] io_tlIn_0_d_bits_data,
  output        io_tlIn_0_d_bits_error,
  output        io_innerCtrl_valid,
  output        io_innerCtrl_bits_resumereq,
  output [9:0]  io_innerCtrl_bits_hartsel
);
  wire [1:0] _T_110;
  wire [23:0] _T_111;
  wire [25:0] _T_112;
  wire [2:0] _T_113;
  wire [1:0] _T_114;
  wire [2:0] _T_115;
  wire [5:0] _T_116;
  wire [31:0] _T_117;
  wire  DMCONTROL_clock;
  wire  DMCONTROL_reset;
  wire [31:0] DMCONTROL_io_d;
  wire [31:0] DMCONTROL_io_q;
  wire  DMCONTROL_io_en;
  wire [31:0] _T_122;
  wire  _T_123;
  wire  _T_124;
  wire [13:0] _T_125;
  wire [9:0] _T_126;
  wire  _T_127;
  wire [1:0] _T_128;
  wire  _T_129;
  wire  _T_130;
  wire  _T_131;
  wire  _T_140;
  wire  _T_141;
  wire [9:0] _T_143;
  wire  _T_147;
  wire  _T_148;
  wire  _T_153;
  wire  _GEN_0;
  wire  _GEN_1;
  wire  _GEN_2;
  wire [1:0] _GEN_3;
  wire  _GEN_4;
  wire [9:0] _GEN_5;
  wire [13:0] _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _T_155;
  wire  _GEN_9;
  wire [9:0] _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [9:0] _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire [1:0] _T_156;
  wire [23:0] _T_157;
  wire [25:0] _T_158;
  wire [2:0] _T_159;
  wire [1:0] _T_160;
  wire [2:0] _T_161;
  wire [5:0] _T_162;
  wire [31:0] _T_163;
  wire  _T_169_bits_index;
  wire  _T_174;
  wire [4:0] _T_175;
  wire [2:0] _T_176;
  wire  _T_203;
  wire  _T_237;
  wire  _T_238;
  wire  _T_239;
  wire  _T_240;
  wire [7:0] _T_244;
  wire [7:0] _T_248;
  wire [7:0] _T_252;
  wire [7:0] _T_256;
  wire [15:0] _T_257;
  wire [15:0] _T_258;
  wire [31:0] _T_259;
  wire [31:0] _T_287;
  wire  _T_289;
  wire  _T_302;
  wire [31:0] _GEN_18;
  wire [1:0] _T_326;
  wire  _T_327;
  wire  _T_333;
  wire  _T_351;
  wire  _T_352;
  wire  _T_355;
  wire  _T_390;
  wire [31:0] _T_432;
  wire  _T_433;
  wire [1:0] _T_434;
  wire  debugInterrupts_clock;
  wire  debugInterrupts_reset;
  wire  debugInterrupts_io_d;
  wire  debugInterrupts_io_q;
  wire  debugInterrupts_io_en;
  wire  _T_469;
  wire  _GEN_19;
  wire  _T_494;
  wire  _T_495;
  wire  _GEN_20;
  wire  _GEN_21;
  AsyncResetRegVec DMCONTROL (
    .clock(DMCONTROL_clock),
    .reset(DMCONTROL_reset),
    .io_d(DMCONTROL_io_d),
    .io_q(DMCONTROL_io_q),
    .io_en(DMCONTROL_io_en)
  );
  AsyncResetRegVec_1 debugInterrupts (
    .clock(debugInterrupts_clock),
    .reset(debugInterrupts_reset),
    .io_d(debugInterrupts_io_d),
    .io_q(debugInterrupts_io_q),
    .io_en(debugInterrupts_io_en)
  );
  assign io_debugInterrupts_0_0 = _T_469;
  assign io_ctrl_ndreset = _T_124;
  assign io_ctrl_dmactive = _T_123;
  assign io_tlIn_0_a_ready = io_tlIn_0_d_ready;
  assign io_tlIn_0_d_valid = io_tlIn_0_a_valid;
  assign io_tlIn_0_d_bits_opcode = {{2'd0}, _T_174};
  assign io_tlIn_0_d_bits_param = 2'h0;
  assign io_tlIn_0_d_bits_size = _T_434;
  assign io_tlIn_0_d_bits_source = _T_433;
  assign io_tlIn_0_d_bits_sink = 1'h0;
  assign io_tlIn_0_d_bits_data = _T_432;
  assign io_tlIn_0_d_bits_error = 1'h0;
  assign io_innerCtrl_valid = _T_302;
  assign io_innerCtrl_bits_resumereq = _T_147;
  assign io_innerCtrl_bits_hartsel = _T_143;
  assign _T_110 = {_GEN_13,_GEN_17};
  assign _T_111 = {_GEN_14,_GEN_6};
  assign _T_112 = {_T_111,_T_110};
  assign _T_113 = {_GEN_3,_GEN_4};
  assign _T_114 = {_GEN_15,_GEN_16};
  assign _T_115 = {_T_114,_GEN_2};
  assign _T_116 = {_T_115,_T_113};
  assign _T_117 = {_T_116,_T_112};
  assign DMCONTROL_clock = clock;
  assign DMCONTROL_reset = reset;
  assign DMCONTROL_io_d = _T_117;
  assign DMCONTROL_io_en = 1'h1;
  assign _T_122 = DMCONTROL_io_q;
  assign _T_123 = _T_122[0];
  assign _T_124 = _T_122[1];
  assign _T_125 = _T_122[15:2];
  assign _T_126 = _T_122[25:16];
  assign _T_127 = _T_122[26];
  assign _T_128 = _T_122[28:27];
  assign _T_129 = _T_122[29];
  assign _T_130 = _T_122[30];
  assign _T_131 = _T_122[31];
  assign _T_140 = _GEN_18[0];
  assign _T_141 = _GEN_18[1];
  assign _T_143 = _GEN_18[25:16];
  assign _T_147 = _GEN_18[30];
  assign _T_148 = _GEN_18[31];
  assign _T_153 = ~ _T_123;
  assign _GEN_0 = _T_153 ? 1'h0 : _T_131;
  assign _GEN_1 = _T_153 ? 1'h0 : _T_130;
  assign _GEN_2 = _T_153 ? 1'h0 : _T_129;
  assign _GEN_3 = _T_153 ? 2'h0 : _T_128;
  assign _GEN_4 = _T_153 ? 1'h0 : _T_127;
  assign _GEN_5 = _T_153 ? 10'h0 : _T_126;
  assign _GEN_6 = _T_153 ? 14'h0 : _T_125;
  assign _GEN_7 = _T_153 ? 1'h0 : _T_124;
  assign _GEN_8 = _T_153 ? 1'h0 : _T_123;
  assign _T_155 = _T_153 == 1'h0;
  assign _GEN_9 = _T_302 ? _T_141 : _GEN_7;
  assign _GEN_10 = _T_302 ? _T_143 : _GEN_5;
  assign _GEN_11 = _T_302 ? _T_148 : _GEN_0;
  assign _GEN_12 = _T_302 ? _T_147 : _GEN_1;
  assign _GEN_13 = _T_155 ? _GEN_9 : _GEN_7;
  assign _GEN_14 = _T_155 ? _GEN_10 : _GEN_5;
  assign _GEN_15 = _T_155 ? _GEN_11 : _GEN_0;
  assign _GEN_16 = _T_155 ? _GEN_12 : _GEN_1;
  assign _GEN_17 = _T_302 ? _T_140 : _GEN_8;
  assign _T_156 = {_T_124,_T_123};
  assign _T_157 = {_T_126,_T_125};
  assign _T_158 = {_T_157,_T_156};
  assign _T_159 = {_T_128,_T_127};
  assign _T_160 = {_T_131,_T_130};
  assign _T_161 = {_T_160,_T_129};
  assign _T_162 = {_T_161,_T_159};
  assign _T_163 = {_T_162,_T_158};
  assign _T_169_bits_index = _T_175[0];
  assign _T_174 = io_tlIn_0_a_bits_opcode == 3'h4;
  assign _T_175 = io_tlIn_0_a_bits_address[6:2];
  assign _T_176 = {io_tlIn_0_a_bits_source,io_tlIn_0_a_bits_size};
  assign _T_203 = _T_169_bits_index == 1'h0;
  assign _T_237 = io_tlIn_0_a_bits_mask[0];
  assign _T_238 = io_tlIn_0_a_bits_mask[1];
  assign _T_239 = io_tlIn_0_a_bits_mask[2];
  assign _T_240 = io_tlIn_0_a_bits_mask[3];
  assign _T_244 = _T_237 ? 8'hff : 8'h0;
  assign _T_248 = _T_238 ? 8'hff : 8'h0;
  assign _T_252 = _T_239 ? 8'hff : 8'h0;
  assign _T_256 = _T_240 ? 8'hff : 8'h0;
  assign _T_257 = {_T_248,_T_244};
  assign _T_258 = {_T_256,_T_252};
  assign _T_259 = {_T_258,_T_257};
  assign _T_287 = ~ _T_259;
  assign _T_289 = _T_287 == 32'h0;
  assign _T_302 = _T_390 & _T_289;
  assign _GEN_18 = _T_302 ? io_tlIn_0_a_bits_data : 32'h0;
  assign _T_326 = 2'h1 << 1'h0;
  assign _T_327 = _T_326[0];
  assign _T_333 = io_tlIn_0_a_valid & io_tlIn_0_d_ready;
  assign _T_351 = _T_174 == 1'h0;
  assign _T_352 = _T_333 & _T_351;
  assign _T_355 = _T_352 & _T_327;
  assign _T_390 = _T_355 & _T_203;
  assign _T_432 = _T_203 ? _T_163 : 32'h0;
  assign _T_433 = _T_176[2];
  assign _T_434 = _T_176[1:0];
  assign debugInterrupts_clock = clock;
  assign debugInterrupts_reset = reset;
  assign debugInterrupts_io_d = _GEN_21;
  assign debugInterrupts_io_en = 1'h1;
  assign _T_469 = debugInterrupts_io_q;
  assign _GEN_19 = _T_153 ? 1'h0 : _T_469;
  assign _T_494 = _T_143 == 10'h0;
  assign _T_495 = _T_302 & _T_494;
  assign _GEN_20 = _T_495 ? _T_148 : _GEN_19;
  assign _GEN_21 = _T_155 ? _GEN_20 : _GEN_19;
endmodule
module AsyncValidSync(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  source_valid_sync_0_clock;
  wire  source_valid_sync_0_reset;
  wire  source_valid_sync_0_io_d;
  wire  source_valid_sync_0_io_q;
  wire  source_valid_sync_0_io_en;
  wire  source_valid_sync_1_clock;
  wire  source_valid_sync_1_reset;
  wire  source_valid_sync_1_io_d;
  wire  source_valid_sync_1_io_q;
  wire  source_valid_sync_1_io_en;
  wire  source_valid_sync_2_clock;
  wire  source_valid_sync_2_reset;
  wire  source_valid_sync_2_io_d;
  wire  source_valid_sync_2_io_q;
  wire  source_valid_sync_2_io_en;
  wire  source_valid_sync_3_clock;
  wire  source_valid_sync_3_reset;
  wire  source_valid_sync_3_io_d;
  wire  source_valid_sync_3_io_q;
  wire  source_valid_sync_3_io_en;
  wire  _T_8;
  AsyncResetRegVec_1 source_valid_sync_0 (
    .clock(source_valid_sync_0_clock),
    .reset(source_valid_sync_0_reset),
    .io_d(source_valid_sync_0_io_d),
    .io_q(source_valid_sync_0_io_q),
    .io_en(source_valid_sync_0_io_en)
  );
  AsyncResetRegVec_1 source_valid_sync_1 (
    .clock(source_valid_sync_1_clock),
    .reset(source_valid_sync_1_reset),
    .io_d(source_valid_sync_1_io_d),
    .io_q(source_valid_sync_1_io_q),
    .io_en(source_valid_sync_1_io_en)
  );
  AsyncResetRegVec_1 source_valid_sync_2 (
    .clock(source_valid_sync_2_clock),
    .reset(source_valid_sync_2_reset),
    .io_d(source_valid_sync_2_io_d),
    .io_q(source_valid_sync_2_io_q),
    .io_en(source_valid_sync_2_io_en)
  );
  AsyncResetRegVec_1 source_valid_sync_3 (
    .clock(source_valid_sync_3_clock),
    .reset(source_valid_sync_3_reset),
    .io_d(source_valid_sync_3_io_d),
    .io_q(source_valid_sync_3_io_q),
    .io_en(source_valid_sync_3_io_en)
  );
  assign io_out = _T_8;
  assign source_valid_sync_0_clock = clock;
  assign source_valid_sync_0_reset = reset;
  assign source_valid_sync_0_io_d = source_valid_sync_1_io_q;
  assign source_valid_sync_0_io_en = 1'h1;
  assign source_valid_sync_1_clock = clock;
  assign source_valid_sync_1_reset = reset;
  assign source_valid_sync_1_io_d = source_valid_sync_2_io_q;
  assign source_valid_sync_1_io_en = 1'h1;
  assign source_valid_sync_2_clock = clock;
  assign source_valid_sync_2_reset = reset;
  assign source_valid_sync_2_io_d = source_valid_sync_3_io_q;
  assign source_valid_sync_2_io_en = 1'h1;
  assign source_valid_sync_3_clock = clock;
  assign source_valid_sync_3_reset = reset;
  assign source_valid_sync_3_io_d = io_in;
  assign source_valid_sync_3_io_en = 1'h1;
  assign _T_8 = source_valid_sync_0_io_q;
endmodule
module AsyncValidSync_1(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sink_extend_sync_0_clock;
  wire  sink_extend_sync_0_reset;
  wire  sink_extend_sync_0_io_d;
  wire  sink_extend_sync_0_io_q;
  wire  sink_extend_sync_0_io_en;
  wire  _T_5;
  AsyncResetRegVec_1 sink_extend_sync_0 (
    .clock(sink_extend_sync_0_clock),
    .reset(sink_extend_sync_0_reset),
    .io_d(sink_extend_sync_0_io_d),
    .io_q(sink_extend_sync_0_io_q),
    .io_en(sink_extend_sync_0_io_en)
  );
  assign io_out = _T_5;
  assign sink_extend_sync_0_clock = clock;
  assign sink_extend_sync_0_reset = reset;
  assign sink_extend_sync_0_io_d = io_in;
  assign sink_extend_sync_0_io_en = 1'h1;
  assign _T_5 = sink_extend_sync_0_io_q;
endmodule
module AsyncValidSync_2(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sink_valid_sync_0_clock;
  wire  sink_valid_sync_0_reset;
  wire  sink_valid_sync_0_io_d;
  wire  sink_valid_sync_0_io_q;
  wire  sink_valid_sync_0_io_en;
  wire  sink_valid_sync_1_clock;
  wire  sink_valid_sync_1_reset;
  wire  sink_valid_sync_1_io_d;
  wire  sink_valid_sync_1_io_q;
  wire  sink_valid_sync_1_io_en;
  wire  sink_valid_sync_2_clock;
  wire  sink_valid_sync_2_reset;
  wire  sink_valid_sync_2_io_d;
  wire  sink_valid_sync_2_io_q;
  wire  sink_valid_sync_2_io_en;
  wire  _T_7;
  AsyncResetRegVec_1 sink_valid_sync_0 (
    .clock(sink_valid_sync_0_clock),
    .reset(sink_valid_sync_0_reset),
    .io_d(sink_valid_sync_0_io_d),
    .io_q(sink_valid_sync_0_io_q),
    .io_en(sink_valid_sync_0_io_en)
  );
  AsyncResetRegVec_1 sink_valid_sync_1 (
    .clock(sink_valid_sync_1_clock),
    .reset(sink_valid_sync_1_reset),
    .io_d(sink_valid_sync_1_io_d),
    .io_q(sink_valid_sync_1_io_q),
    .io_en(sink_valid_sync_1_io_en)
  );
  AsyncResetRegVec_1 sink_valid_sync_2 (
    .clock(sink_valid_sync_2_clock),
    .reset(sink_valid_sync_2_reset),
    .io_d(sink_valid_sync_2_io_d),
    .io_q(sink_valid_sync_2_io_q),
    .io_en(sink_valid_sync_2_io_en)
  );
  assign io_out = _T_7;
  assign sink_valid_sync_0_clock = clock;
  assign sink_valid_sync_0_reset = reset;
  assign sink_valid_sync_0_io_d = sink_valid_sync_1_io_q;
  assign sink_valid_sync_0_io_en = 1'h1;
  assign sink_valid_sync_1_clock = clock;
  assign sink_valid_sync_1_reset = reset;
  assign sink_valid_sync_1_io_d = sink_valid_sync_2_io_q;
  assign sink_valid_sync_1_io_en = 1'h1;
  assign sink_valid_sync_2_clock = clock;
  assign sink_valid_sync_2_reset = reset;
  assign sink_valid_sync_2_io_d = io_in;
  assign sink_valid_sync_2_io_en = 1'h1;
  assign _T_7 = sink_valid_sync_0_io_q;
endmodule
module AsyncQueueSource(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_size,
  input         io_enq_bits_source,
  input  [8:0]  io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_ridx,
  output        io_widx,
  output [2:0]  io_mem_0_opcode,
  output [1:0]  io_mem_0_size,
  output        io_mem_0_source,
  output [8:0]  io_mem_0_address,
  output [3:0]  io_mem_0_mask,
  output [31:0] io_mem_0_data,
  input         io_sink_reset_n,
  input         io_ridx_valid,
  output        io_widx_valid
);
  wire  sink_ready;
  reg [2:0] mem_0_opcode;
  reg [31:0] _RAND_0;
  reg [1:0] mem_0_size;
  reg [31:0] _RAND_1;
  reg  mem_0_source;
  reg [31:0] _RAND_2;
  reg [8:0] mem_0_address;
  reg [31:0] _RAND_3;
  reg [3:0] mem_0_mask;
  reg [31:0] _RAND_4;
  reg [31:0] mem_0_data;
  reg [31:0] _RAND_5;
  wire  _T_26;
  wire  _T_28;
  wire  widx_bin_clock;
  wire  widx_bin_reset;
  wire  widx_bin_io_d;
  wire  widx_bin_io_q;
  wire  widx_bin_io_en;
  wire [1:0] _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_37;
  wire  widx;
  wire  ridx_gray_sync_0_clock;
  wire  ridx_gray_sync_0_reset;
  wire  ridx_gray_sync_0_io_d;
  wire  ridx_gray_sync_0_io_q;
  wire  ridx_gray_sync_0_io_en;
  wire  ridx_gray_sync_1_clock;
  wire  ridx_gray_sync_1_reset;
  wire  ridx_gray_sync_1_io_d;
  wire  ridx_gray_sync_1_io_q;
  wire  ridx_gray_sync_1_io_en;
  wire  ridx_gray_sync_2_clock;
  wire  ridx_gray_sync_2_reset;
  wire  ridx_gray_sync_2_io_d;
  wire  ridx_gray_sync_2_io_q;
  wire  ridx_gray_sync_2_io_en;
  wire  _T_42;
  wire  _T_43;
  wire  ready;
  wire [2:0] _GEN_0;
  wire [1:0] _GEN_2;
  wire  _GEN_3;
  wire [8:0] _GEN_4;
  wire [3:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire  ready_reg_clock;
  wire  ready_reg_reset;
  wire  ready_reg_io_d;
  wire  ready_reg_io_q;
  wire  ready_reg_io_en;
  wire  ready_reg_1;
  wire  _T_48;
  wire  widx_gray_clock;
  wire  widx_gray_reset;
  wire  widx_gray_io_d;
  wire  widx_gray_io_q;
  wire  widx_gray_io_en;
  wire  AsyncValidSync_clock;
  wire  AsyncValidSync_reset;
  wire  AsyncValidSync_io_in;
  wire  AsyncValidSync_io_out;
  wire  AsyncValidSync_1_clock;
  wire  AsyncValidSync_1_reset;
  wire  AsyncValidSync_1_io_in;
  wire  AsyncValidSync_1_io_out;
  wire  AsyncValidSync_2_clock;
  wire  AsyncValidSync_2_reset;
  wire  AsyncValidSync_2_io_in;
  wire  AsyncValidSync_2_io_out;
  wire  _T_52;
  wire  _T_53;
  AsyncResetRegVec_1 widx_bin (
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_0 (
    .clock(ridx_gray_sync_0_clock),
    .reset(ridx_gray_sync_0_reset),
    .io_d(ridx_gray_sync_0_io_d),
    .io_q(ridx_gray_sync_0_io_q),
    .io_en(ridx_gray_sync_0_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_1 (
    .clock(ridx_gray_sync_1_clock),
    .reset(ridx_gray_sync_1_reset),
    .io_d(ridx_gray_sync_1_io_d),
    .io_q(ridx_gray_sync_1_io_q),
    .io_en(ridx_gray_sync_1_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_2 (
    .clock(ridx_gray_sync_2_clock),
    .reset(ridx_gray_sync_2_reset),
    .io_d(ridx_gray_sync_2_io_d),
    .io_q(ridx_gray_sync_2_io_q),
    .io_en(ridx_gray_sync_2_io_en)
  );
  AsyncResetRegVec_1 ready_reg (
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_1 widx_gray (
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync (
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 (
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 (
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign io_enq_ready = _T_48;
  assign io_widx = widx_gray_io_q;
  assign io_mem_0_opcode = mem_0_opcode;
  assign io_mem_0_size = mem_0_size;
  assign io_mem_0_source = mem_0_source;
  assign io_mem_0_address = mem_0_address;
  assign io_mem_0_mask = mem_0_mask;
  assign io_mem_0_data = mem_0_data;
  assign io_widx_valid = AsyncValidSync_io_out;
  assign sink_ready = AsyncValidSync_2_io_out;
  assign _T_26 = io_enq_ready & io_enq_valid;
  assign _T_28 = sink_ready == 1'h0;
  assign widx_bin_clock = clock;
  assign widx_bin_reset = reset;
  assign widx_bin_io_d = _T_35;
  assign widx_bin_io_en = 1'h1;
  assign _T_33 = widx_bin_io_q + _T_26;
  assign _T_34 = _T_33[0:0];
  assign _T_35 = _T_28 ? 1'h0 : _T_34;
  assign _T_37 = _T_35 >> 1'h1;
  assign widx = _T_35 ^ _T_37;
  assign ridx_gray_sync_0_clock = clock;
  assign ridx_gray_sync_0_reset = reset;
  assign ridx_gray_sync_0_io_d = ridx_gray_sync_1_io_q;
  assign ridx_gray_sync_0_io_en = 1'h1;
  assign ridx_gray_sync_1_clock = clock;
  assign ridx_gray_sync_1_reset = reset;
  assign ridx_gray_sync_1_io_d = ridx_gray_sync_2_io_q;
  assign ridx_gray_sync_1_io_en = 1'h1;
  assign ridx_gray_sync_2_clock = clock;
  assign ridx_gray_sync_2_reset = reset;
  assign ridx_gray_sync_2_io_d = io_ridx;
  assign ridx_gray_sync_2_io_en = 1'h1;
  assign _T_42 = ridx_gray_sync_0_io_q ^ 1'h1;
  assign _T_43 = widx != _T_42;
  assign ready = sink_ready & _T_43;
  assign _GEN_0 = _T_26 ? io_enq_bits_opcode : mem_0_opcode;
  assign _GEN_2 = _T_26 ? io_enq_bits_size : mem_0_size;
  assign _GEN_3 = _T_26 ? io_enq_bits_source : mem_0_source;
  assign _GEN_4 = _T_26 ? io_enq_bits_address : mem_0_address;
  assign _GEN_5 = _T_26 ? io_enq_bits_mask : mem_0_mask;
  assign _GEN_6 = _T_26 ? io_enq_bits_data : mem_0_data;
  assign ready_reg_clock = clock;
  assign ready_reg_reset = reset;
  assign ready_reg_io_d = ready;
  assign ready_reg_io_en = 1'h1;
  assign ready_reg_1 = ready_reg_io_q;
  assign _T_48 = ready_reg_1 & sink_ready;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = widx;
  assign widx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_53;
  assign AsyncValidSync_io_in = 1'h1;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_53;
  assign AsyncValidSync_1_io_in = io_ridx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign _T_52 = io_sink_reset_n == 1'h0;
  assign _T_53 = reset | _T_52;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  mem_0_opcode = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0_size = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem_0_source = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_0_address = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  mem_0_mask = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_0_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_26) begin
      mem_0_opcode <= io_enq_bits_opcode;
    end
    if (_T_26) begin
      mem_0_size <= io_enq_bits_size;
    end
    if (_T_26) begin
      mem_0_source <= io_enq_bits_source;
    end
    if (_T_26) begin
      mem_0_address <= io_enq_bits_address;
    end
    if (_T_26) begin
      mem_0_mask <= io_enq_bits_mask;
    end
    if (_T_26) begin
      mem_0_data <= io_enq_bits_data;
    end
  end
endmodule
module AsyncValidSync_3(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sink_valid_sync_0_clock;
  wire  sink_valid_sync_0_reset;
  wire  sink_valid_sync_0_io_d;
  wire  sink_valid_sync_0_io_q;
  wire  sink_valid_sync_0_io_en;
  wire  sink_valid_sync_1_clock;
  wire  sink_valid_sync_1_reset;
  wire  sink_valid_sync_1_io_d;
  wire  sink_valid_sync_1_io_q;
  wire  sink_valid_sync_1_io_en;
  wire  sink_valid_sync_2_clock;
  wire  sink_valid_sync_2_reset;
  wire  sink_valid_sync_2_io_d;
  wire  sink_valid_sync_2_io_q;
  wire  sink_valid_sync_2_io_en;
  wire  sink_valid_sync_3_clock;
  wire  sink_valid_sync_3_reset;
  wire  sink_valid_sync_3_io_d;
  wire  sink_valid_sync_3_io_q;
  wire  sink_valid_sync_3_io_en;
  wire  _T_8;
  AsyncResetRegVec_1 sink_valid_sync_0 (
    .clock(sink_valid_sync_0_clock),
    .reset(sink_valid_sync_0_reset),
    .io_d(sink_valid_sync_0_io_d),
    .io_q(sink_valid_sync_0_io_q),
    .io_en(sink_valid_sync_0_io_en)
  );
  AsyncResetRegVec_1 sink_valid_sync_1 (
    .clock(sink_valid_sync_1_clock),
    .reset(sink_valid_sync_1_reset),
    .io_d(sink_valid_sync_1_io_d),
    .io_q(sink_valid_sync_1_io_q),
    .io_en(sink_valid_sync_1_io_en)
  );
  AsyncResetRegVec_1 sink_valid_sync_2 (
    .clock(sink_valid_sync_2_clock),
    .reset(sink_valid_sync_2_reset),
    .io_d(sink_valid_sync_2_io_d),
    .io_q(sink_valid_sync_2_io_q),
    .io_en(sink_valid_sync_2_io_en)
  );
  AsyncResetRegVec_1 sink_valid_sync_3 (
    .clock(sink_valid_sync_3_clock),
    .reset(sink_valid_sync_3_reset),
    .io_d(sink_valid_sync_3_io_d),
    .io_q(sink_valid_sync_3_io_q),
    .io_en(sink_valid_sync_3_io_en)
  );
  assign io_out = _T_8;
  assign sink_valid_sync_0_clock = clock;
  assign sink_valid_sync_0_reset = reset;
  assign sink_valid_sync_0_io_d = sink_valid_sync_1_io_q;
  assign sink_valid_sync_0_io_en = 1'h1;
  assign sink_valid_sync_1_clock = clock;
  assign sink_valid_sync_1_reset = reset;
  assign sink_valid_sync_1_io_d = sink_valid_sync_2_io_q;
  assign sink_valid_sync_1_io_en = 1'h1;
  assign sink_valid_sync_2_clock = clock;
  assign sink_valid_sync_2_reset = reset;
  assign sink_valid_sync_2_io_d = sink_valid_sync_3_io_q;
  assign sink_valid_sync_2_io_en = 1'h1;
  assign sink_valid_sync_3_clock = clock;
  assign sink_valid_sync_3_reset = reset;
  assign sink_valid_sync_3_io_d = io_in;
  assign sink_valid_sync_3_io_en = 1'h1;
  assign _T_8 = sink_valid_sync_0_io_q;
endmodule
module AsyncValidSync_4(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  source_extend_sync_0_clock;
  wire  source_extend_sync_0_reset;
  wire  source_extend_sync_0_io_d;
  wire  source_extend_sync_0_io_q;
  wire  source_extend_sync_0_io_en;
  wire  _T_5;
  AsyncResetRegVec_1 source_extend_sync_0 (
    .clock(source_extend_sync_0_clock),
    .reset(source_extend_sync_0_reset),
    .io_d(source_extend_sync_0_io_d),
    .io_q(source_extend_sync_0_io_q),
    .io_en(source_extend_sync_0_io_en)
  );
  assign io_out = _T_5;
  assign source_extend_sync_0_clock = clock;
  assign source_extend_sync_0_reset = reset;
  assign source_extend_sync_0_io_d = io_in;
  assign source_extend_sync_0_io_en = 1'h1;
  assign _T_5 = source_extend_sync_0_io_q;
endmodule
module AsyncValidSync_5(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  source_valid_sync_0_clock;
  wire  source_valid_sync_0_reset;
  wire  source_valid_sync_0_io_d;
  wire  source_valid_sync_0_io_q;
  wire  source_valid_sync_0_io_en;
  wire  source_valid_sync_1_clock;
  wire  source_valid_sync_1_reset;
  wire  source_valid_sync_1_io_d;
  wire  source_valid_sync_1_io_q;
  wire  source_valid_sync_1_io_en;
  wire  source_valid_sync_2_clock;
  wire  source_valid_sync_2_reset;
  wire  source_valid_sync_2_io_d;
  wire  source_valid_sync_2_io_q;
  wire  source_valid_sync_2_io_en;
  wire  _T_7;
  AsyncResetRegVec_1 source_valid_sync_0 (
    .clock(source_valid_sync_0_clock),
    .reset(source_valid_sync_0_reset),
    .io_d(source_valid_sync_0_io_d),
    .io_q(source_valid_sync_0_io_q),
    .io_en(source_valid_sync_0_io_en)
  );
  AsyncResetRegVec_1 source_valid_sync_1 (
    .clock(source_valid_sync_1_clock),
    .reset(source_valid_sync_1_reset),
    .io_d(source_valid_sync_1_io_d),
    .io_q(source_valid_sync_1_io_q),
    .io_en(source_valid_sync_1_io_en)
  );
  AsyncResetRegVec_1 source_valid_sync_2 (
    .clock(source_valid_sync_2_clock),
    .reset(source_valid_sync_2_reset),
    .io_d(source_valid_sync_2_io_d),
    .io_q(source_valid_sync_2_io_q),
    .io_en(source_valid_sync_2_io_en)
  );
  assign io_out = _T_7;
  assign source_valid_sync_0_clock = clock;
  assign source_valid_sync_0_reset = reset;
  assign source_valid_sync_0_io_d = source_valid_sync_1_io_q;
  assign source_valid_sync_0_io_en = 1'h1;
  assign source_valid_sync_1_clock = clock;
  assign source_valid_sync_1_reset = reset;
  assign source_valid_sync_1_io_d = source_valid_sync_2_io_q;
  assign source_valid_sync_1_io_en = 1'h1;
  assign source_valid_sync_2_clock = clock;
  assign source_valid_sync_2_reset = reset;
  assign source_valid_sync_2_io_d = io_in;
  assign source_valid_sync_2_io_en = 1'h1;
  assign _T_7 = source_valid_sync_0_io_q;
endmodule
module AsyncQueueSink(
  input         clock,
  input         reset,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [1:0]  io_deq_bits_size,
  output        io_deq_bits_source,
  output        io_deq_bits_sink,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_error,
  output        io_ridx,
  input         io_widx,
  input  [2:0]  io_mem_0_opcode,
  input  [1:0]  io_mem_0_param,
  input  [1:0]  io_mem_0_size,
  input         io_mem_0_source,
  input         io_mem_0_sink,
  input  [31:0] io_mem_0_data,
  input         io_mem_0_error,
  input         io_source_reset_n,
  output        io_ridx_valid,
  input         io_widx_valid
);
  wire  source_ready;
  wire  _T_17;
  wire  _T_19;
  wire  ridx_bin_clock;
  wire  ridx_bin_reset;
  wire  ridx_bin_io_d;
  wire  ridx_bin_io_q;
  wire  ridx_bin_io_en;
  wire [1:0] _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_28;
  wire  ridx;
  wire  widx_gray_sync_0_clock;
  wire  widx_gray_sync_0_reset;
  wire  widx_gray_sync_0_io_d;
  wire  widx_gray_sync_0_io_q;
  wire  widx_gray_sync_0_io_en;
  wire  widx_gray_sync_1_clock;
  wire  widx_gray_sync_1_reset;
  wire  widx_gray_sync_1_io_d;
  wire  widx_gray_sync_1_io_q;
  wire  widx_gray_sync_1_io_en;
  wire  widx_gray_sync_2_clock;
  wire  widx_gray_sync_2_reset;
  wire  widx_gray_sync_2_io_d;
  wire  widx_gray_sync_2_io_q;
  wire  widx_gray_sync_2_io_en;
  wire  _T_32;
  wire  valid;
  reg [2:0] _T_36_opcode;
  reg [31:0] _RAND_0;
  reg [1:0] _T_36_param;
  reg [31:0] _RAND_1;
  reg [1:0] _T_36_size;
  reg [31:0] _RAND_2;
  reg  _T_36_source;
  reg [31:0] _RAND_3;
  reg  _T_36_sink;
  reg [31:0] _RAND_4;
  reg [31:0] _T_36_data;
  reg [31:0] _RAND_5;
  reg  _T_36_error;
  reg [31:0] _RAND_6;
  wire [2:0] _GEN_0;
  wire [1:0] _GEN_1;
  wire [1:0] _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [31:0] _GEN_5;
  wire  _GEN_6;
  wire  valid_reg_clock;
  wire  valid_reg_reset;
  wire  valid_reg_io_d;
  wire  valid_reg_io_q;
  wire  valid_reg_io_en;
  wire  valid_reg_1;
  wire  _T_38;
  wire  ridx_gray_clock;
  wire  ridx_gray_reset;
  wire  ridx_gray_io_d;
  wire  ridx_gray_io_q;
  wire  ridx_gray_io_en;
  wire  AsyncValidSync_clock;
  wire  AsyncValidSync_reset;
  wire  AsyncValidSync_io_in;
  wire  AsyncValidSync_io_out;
  wire  AsyncValidSync_1_clock;
  wire  AsyncValidSync_1_reset;
  wire  AsyncValidSync_1_io_in;
  wire  AsyncValidSync_1_io_out;
  wire  AsyncValidSync_2_clock;
  wire  AsyncValidSync_2_reset;
  wire  AsyncValidSync_2_io_in;
  wire  AsyncValidSync_2_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  _T_60;
  wire  AsyncResetRegVec_clock;
  wire  AsyncResetRegVec_reset;
  wire  AsyncResetRegVec_io_d;
  wire  AsyncResetRegVec_io_q;
  wire  AsyncResetRegVec_io_en;
  AsyncResetRegVec_1 ridx_bin (
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_0 (
    .clock(widx_gray_sync_0_clock),
    .reset(widx_gray_sync_0_reset),
    .io_d(widx_gray_sync_0_io_d),
    .io_q(widx_gray_sync_0_io_q),
    .io_en(widx_gray_sync_0_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_1 (
    .clock(widx_gray_sync_1_clock),
    .reset(widx_gray_sync_1_reset),
    .io_d(widx_gray_sync_1_io_d),
    .io_q(widx_gray_sync_1_io_q),
    .io_en(widx_gray_sync_1_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_2 (
    .clock(widx_gray_sync_2_clock),
    .reset(widx_gray_sync_2_reset),
    .io_d(widx_gray_sync_2_io_d),
    .io_q(widx_gray_sync_2_io_q),
    .io_en(widx_gray_sync_2_io_en)
  );
  AsyncResetRegVec_1 valid_reg (
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_1 ridx_gray (
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync_3 AsyncValidSync (
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_4 AsyncValidSync_1 (
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_5 AsyncValidSync_2 (
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_1 AsyncResetRegVec (
    .clock(AsyncResetRegVec_clock),
    .reset(AsyncResetRegVec_reset),
    .io_d(AsyncResetRegVec_io_d),
    .io_q(AsyncResetRegVec_io_q),
    .io_en(AsyncResetRegVec_io_en)
  );
  assign io_deq_valid = _T_38;
  assign io_deq_bits_opcode = _T_36_opcode;
  assign io_deq_bits_param = _T_36_param;
  assign io_deq_bits_size = _T_36_size;
  assign io_deq_bits_source = _T_36_source;
  assign io_deq_bits_sink = _T_36_sink;
  assign io_deq_bits_data = _T_36_data;
  assign io_deq_bits_error = _T_36_error;
  assign io_ridx = ridx_gray_io_q;
  assign io_ridx_valid = AsyncValidSync_io_out;
  assign source_ready = AsyncValidSync_2_io_out;
  assign _T_17 = io_deq_ready & io_deq_valid;
  assign _T_19 = source_ready == 1'h0;
  assign ridx_bin_clock = clock;
  assign ridx_bin_reset = reset;
  assign ridx_bin_io_d = _T_26;
  assign ridx_bin_io_en = 1'h1;
  assign _T_24 = ridx_bin_io_q + _T_17;
  assign _T_25 = _T_24[0:0];
  assign _T_26 = _T_19 ? 1'h0 : _T_25;
  assign _T_28 = _T_26 >> 1'h1;
  assign ridx = _T_26 ^ _T_28;
  assign widx_gray_sync_0_clock = clock;
  assign widx_gray_sync_0_reset = reset;
  assign widx_gray_sync_0_io_d = widx_gray_sync_1_io_q;
  assign widx_gray_sync_0_io_en = 1'h1;
  assign widx_gray_sync_1_clock = clock;
  assign widx_gray_sync_1_reset = reset;
  assign widx_gray_sync_1_io_d = widx_gray_sync_2_io_q;
  assign widx_gray_sync_1_io_en = 1'h1;
  assign widx_gray_sync_2_clock = clock;
  assign widx_gray_sync_2_reset = reset;
  assign widx_gray_sync_2_io_d = io_widx;
  assign widx_gray_sync_2_io_en = 1'h1;
  assign _T_32 = ridx != widx_gray_sync_0_io_q;
  assign valid = source_ready & _T_32;
  assign _GEN_0 = valid ? io_mem_0_opcode : _T_36_opcode;
  assign _GEN_1 = valid ? io_mem_0_param : _T_36_param;
  assign _GEN_2 = valid ? io_mem_0_size : _T_36_size;
  assign _GEN_3 = valid ? io_mem_0_source : _T_36_source;
  assign _GEN_4 = valid ? io_mem_0_sink : _T_36_sink;
  assign _GEN_5 = valid ? io_mem_0_data : _T_36_data;
  assign _GEN_6 = valid ? io_mem_0_error : _T_36_error;
  assign valid_reg_clock = clock;
  assign valid_reg_reset = reset;
  assign valid_reg_io_d = valid;
  assign valid_reg_io_en = 1'h1;
  assign valid_reg_1 = valid_reg_io_q;
  assign _T_38 = valid_reg_1 & source_ready;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = ridx;
  assign ridx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_43;
  assign AsyncValidSync_io_in = 1'h1;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_43;
  assign AsyncValidSync_1_io_in = io_widx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign _T_42 = io_source_reset_n == 1'h0;
  assign _T_43 = reset | _T_42;
  assign _T_60 = io_widx == io_ridx;
  assign AsyncResetRegVec_clock = clock;
  assign AsyncResetRegVec_reset = reset;
  assign AsyncResetRegVec_io_d = _T_60;
  assign AsyncResetRegVec_io_en = 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_36_opcode = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_36_param = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_36_size = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_36_source = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_36_sink = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_36_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_36_error = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (valid) begin
      _T_36_opcode <= io_mem_0_opcode;
    end
    if (valid) begin
      _T_36_param <= io_mem_0_param;
    end
    if (valid) begin
      _T_36_size <= io_mem_0_size;
    end
    if (valid) begin
      _T_36_source <= io_mem_0_source;
    end
    if (valid) begin
      _T_36_sink <= io_mem_0_sink;
    end
    if (valid) begin
      _T_36_data <= io_mem_0_data;
    end
    if (valid) begin
      _T_36_error <= io_mem_0_error;
    end
  end
endmodule
module TLAsyncCrossingSource_dmInner(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [1:0]  io_in_0_a_bits_size,
  input         io_in_0_a_bits_source,
  input  [8:0]  io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [1:0]  io_in_0_d_bits_size,
  output        io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  output [2:0]  io_out_0_a_mem_0_opcode,
  output [1:0]  io_out_0_a_mem_0_size,
  output        io_out_0_a_mem_0_source,
  output [8:0]  io_out_0_a_mem_0_address,
  output [3:0]  io_out_0_a_mem_0_mask,
  output [31:0] io_out_0_a_mem_0_data,
  input         io_out_0_a_ridx,
  output        io_out_0_a_widx,
  input         io_out_0_a_ridx_valid,
  output        io_out_0_a_widx_valid,
  output        io_out_0_a_source_reset_n,
  input         io_out_0_a_sink_reset_n,
  input  [2:0]  io_out_0_d_mem_0_opcode,
  input  [1:0]  io_out_0_d_mem_0_param,
  input  [1:0]  io_out_0_d_mem_0_size,
  input         io_out_0_d_mem_0_source,
  input         io_out_0_d_mem_0_sink,
  input  [31:0] io_out_0_d_mem_0_data,
  input         io_out_0_d_mem_0_error,
  output        io_out_0_d_ridx,
  input         io_out_0_d_widx,
  output        io_out_0_d_ridx_valid,
  input         io_out_0_d_widx_valid,
  input         io_out_0_d_source_reset_n,
  output        io_out_0_d_sink_reset_n
);
  wire  AsyncQueueSource_clock;
  wire  AsyncQueueSource_reset;
  wire  AsyncQueueSource_io_enq_ready;
  wire  AsyncQueueSource_io_enq_valid;
  wire [2:0] AsyncQueueSource_io_enq_bits_opcode;
  wire [1:0] AsyncQueueSource_io_enq_bits_size;
  wire  AsyncQueueSource_io_enq_bits_source;
  wire [8:0] AsyncQueueSource_io_enq_bits_address;
  wire [3:0] AsyncQueueSource_io_enq_bits_mask;
  wire [31:0] AsyncQueueSource_io_enq_bits_data;
  wire  AsyncQueueSource_io_ridx;
  wire  AsyncQueueSource_io_widx;
  wire [2:0] AsyncQueueSource_io_mem_0_opcode;
  wire [1:0] AsyncQueueSource_io_mem_0_size;
  wire  AsyncQueueSource_io_mem_0_source;
  wire [8:0] AsyncQueueSource_io_mem_0_address;
  wire [3:0] AsyncQueueSource_io_mem_0_mask;
  wire [31:0] AsyncQueueSource_io_mem_0_data;
  wire  AsyncQueueSource_io_sink_reset_n;
  wire  AsyncQueueSource_io_ridx_valid;
  wire  AsyncQueueSource_io_widx_valid;
  wire [2:0] _T_102_mem_0_opcode;
  wire [1:0] _T_102_mem_0_size;
  wire  _T_102_mem_0_source;
  wire [8:0] _T_102_mem_0_address;
  wire [3:0] _T_102_mem_0_mask;
  wire [31:0] _T_102_mem_0_data;
  wire  _T_102_widx;
  wire  _T_102_widx_valid;
  wire  _T_108;
  wire  AsyncQueueSink_clock;
  wire  AsyncQueueSink_reset;
  wire  AsyncQueueSink_io_deq_ready;
  wire  AsyncQueueSink_io_deq_valid;
  wire [2:0] AsyncQueueSink_io_deq_bits_opcode;
  wire [1:0] AsyncQueueSink_io_deq_bits_param;
  wire [1:0] AsyncQueueSink_io_deq_bits_size;
  wire  AsyncQueueSink_io_deq_bits_source;
  wire  AsyncQueueSink_io_deq_bits_sink;
  wire [31:0] AsyncQueueSink_io_deq_bits_data;
  wire  AsyncQueueSink_io_deq_bits_error;
  wire  AsyncQueueSink_io_ridx;
  wire  AsyncQueueSink_io_widx;
  wire [2:0] AsyncQueueSink_io_mem_0_opcode;
  wire [1:0] AsyncQueueSink_io_mem_0_param;
  wire [1:0] AsyncQueueSink_io_mem_0_size;
  wire  AsyncQueueSink_io_mem_0_source;
  wire  AsyncQueueSink_io_mem_0_sink;
  wire [31:0] AsyncQueueSink_io_mem_0_data;
  wire  AsyncQueueSink_io_mem_0_error;
  wire  AsyncQueueSink_io_source_reset_n;
  wire  AsyncQueueSink_io_ridx_valid;
  wire  AsyncQueueSink_io_widx_valid;
  wire  _T_110;
  wire  _T_115_valid;
  wire [2:0] _T_115_bits_opcode;
  wire [1:0] _T_115_bits_param;
  wire [1:0] _T_115_bits_size;
  wire  _T_115_bits_source;
  wire  _T_115_bits_sink;
  wire [31:0] _T_115_bits_data;
  wire  _T_115_bits_error;
  AsyncQueueSource AsyncQueueSource (
    .clock(AsyncQueueSource_clock),
    .reset(AsyncQueueSource_reset),
    .io_enq_ready(AsyncQueueSource_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_io_enq_valid),
    .io_enq_bits_opcode(AsyncQueueSource_io_enq_bits_opcode),
    .io_enq_bits_size(AsyncQueueSource_io_enq_bits_size),
    .io_enq_bits_source(AsyncQueueSource_io_enq_bits_source),
    .io_enq_bits_address(AsyncQueueSource_io_enq_bits_address),
    .io_enq_bits_mask(AsyncQueueSource_io_enq_bits_mask),
    .io_enq_bits_data(AsyncQueueSource_io_enq_bits_data),
    .io_ridx(AsyncQueueSource_io_ridx),
    .io_widx(AsyncQueueSource_io_widx),
    .io_mem_0_opcode(AsyncQueueSource_io_mem_0_opcode),
    .io_mem_0_size(AsyncQueueSource_io_mem_0_size),
    .io_mem_0_source(AsyncQueueSource_io_mem_0_source),
    .io_mem_0_address(AsyncQueueSource_io_mem_0_address),
    .io_mem_0_mask(AsyncQueueSource_io_mem_0_mask),
    .io_mem_0_data(AsyncQueueSource_io_mem_0_data),
    .io_sink_reset_n(AsyncQueueSource_io_sink_reset_n),
    .io_ridx_valid(AsyncQueueSource_io_ridx_valid),
    .io_widx_valid(AsyncQueueSource_io_widx_valid)
  );
  AsyncQueueSink AsyncQueueSink (
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits_opcode(AsyncQueueSink_io_deq_bits_opcode),
    .io_deq_bits_param(AsyncQueueSink_io_deq_bits_param),
    .io_deq_bits_size(AsyncQueueSink_io_deq_bits_size),
    .io_deq_bits_source(AsyncQueueSink_io_deq_bits_source),
    .io_deq_bits_sink(AsyncQueueSink_io_deq_bits_sink),
    .io_deq_bits_data(AsyncQueueSink_io_deq_bits_data),
    .io_deq_bits_error(AsyncQueueSink_io_deq_bits_error),
    .io_ridx(AsyncQueueSink_io_ridx),
    .io_widx(AsyncQueueSink_io_widx),
    .io_mem_0_opcode(AsyncQueueSink_io_mem_0_opcode),
    .io_mem_0_param(AsyncQueueSink_io_mem_0_param),
    .io_mem_0_size(AsyncQueueSink_io_mem_0_size),
    .io_mem_0_source(AsyncQueueSink_io_mem_0_source),
    .io_mem_0_sink(AsyncQueueSink_io_mem_0_sink),
    .io_mem_0_data(AsyncQueueSink_io_mem_0_data),
    .io_mem_0_error(AsyncQueueSink_io_mem_0_error),
    .io_source_reset_n(AsyncQueueSink_io_source_reset_n),
    .io_ridx_valid(AsyncQueueSink_io_ridx_valid),
    .io_widx_valid(AsyncQueueSink_io_widx_valid)
  );
  assign io_in_0_a_ready = AsyncQueueSource_io_enq_ready;
  assign io_in_0_d_valid = _T_115_valid;
  assign io_in_0_d_bits_opcode = _T_115_bits_opcode;
  assign io_in_0_d_bits_param = _T_115_bits_param;
  assign io_in_0_d_bits_size = _T_115_bits_size;
  assign io_in_0_d_bits_source = _T_115_bits_source;
  assign io_in_0_d_bits_sink = _T_115_bits_sink;
  assign io_in_0_d_bits_data = _T_115_bits_data;
  assign io_in_0_d_bits_error = _T_115_bits_error;
  assign io_out_0_a_mem_0_opcode = _T_102_mem_0_opcode;
  assign io_out_0_a_mem_0_size = _T_102_mem_0_size;
  assign io_out_0_a_mem_0_source = _T_102_mem_0_source;
  assign io_out_0_a_mem_0_address = _T_102_mem_0_address;
  assign io_out_0_a_mem_0_mask = _T_102_mem_0_mask;
  assign io_out_0_a_mem_0_data = _T_102_mem_0_data;
  assign io_out_0_a_widx = _T_102_widx;
  assign io_out_0_a_widx_valid = _T_102_widx_valid;
  assign io_out_0_a_source_reset_n = _T_108;
  assign io_out_0_d_ridx = AsyncQueueSink_io_ridx;
  assign io_out_0_d_ridx_valid = AsyncQueueSink_io_ridx_valid;
  assign io_out_0_d_sink_reset_n = _T_110;
  assign AsyncQueueSource_clock = clock;
  assign AsyncQueueSource_reset = reset;
  assign AsyncQueueSource_io_enq_valid = io_in_0_a_valid;
  assign AsyncQueueSource_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign AsyncQueueSource_io_enq_bits_size = io_in_0_a_bits_size;
  assign AsyncQueueSource_io_enq_bits_source = io_in_0_a_bits_source;
  assign AsyncQueueSource_io_enq_bits_address = io_in_0_a_bits_address;
  assign AsyncQueueSource_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign AsyncQueueSource_io_enq_bits_data = io_in_0_a_bits_data;
  assign AsyncQueueSource_io_ridx = io_out_0_a_ridx;
  assign AsyncQueueSource_io_sink_reset_n = io_out_0_a_sink_reset_n;
  assign AsyncQueueSource_io_ridx_valid = io_out_0_a_ridx_valid;
  assign _T_102_mem_0_opcode = AsyncQueueSource_io_mem_0_opcode;
  assign _T_102_mem_0_size = AsyncQueueSource_io_mem_0_size;
  assign _T_102_mem_0_source = AsyncQueueSource_io_mem_0_source;
  assign _T_102_mem_0_address = AsyncQueueSource_io_mem_0_address;
  assign _T_102_mem_0_mask = AsyncQueueSource_io_mem_0_mask;
  assign _T_102_mem_0_data = AsyncQueueSource_io_mem_0_data;
  assign _T_102_widx = AsyncQueueSource_io_widx;
  assign _T_102_widx_valid = AsyncQueueSource_io_widx_valid;
  assign _T_108 = AsyncQueueSource_reset == 1'h0;
  assign AsyncQueueSink_clock = clock;
  assign AsyncQueueSink_reset = reset;
  assign AsyncQueueSink_io_deq_ready = io_in_0_d_ready;
  assign AsyncQueueSink_io_widx = io_out_0_d_widx;
  assign AsyncQueueSink_io_mem_0_opcode = io_out_0_d_mem_0_opcode;
  assign AsyncQueueSink_io_mem_0_param = io_out_0_d_mem_0_param;
  assign AsyncQueueSink_io_mem_0_size = io_out_0_d_mem_0_size;
  assign AsyncQueueSink_io_mem_0_source = io_out_0_d_mem_0_source;
  assign AsyncQueueSink_io_mem_0_sink = io_out_0_d_mem_0_sink;
  assign AsyncQueueSink_io_mem_0_data = io_out_0_d_mem_0_data;
  assign AsyncQueueSink_io_mem_0_error = io_out_0_d_mem_0_error;
  assign AsyncQueueSink_io_source_reset_n = io_out_0_d_source_reset_n;
  assign AsyncQueueSink_io_widx_valid = io_out_0_d_widx_valid;
  assign _T_110 = AsyncQueueSink_reset == 1'h0;
  assign _T_115_valid = AsyncQueueSink_io_deq_valid;
  assign _T_115_bits_opcode = AsyncQueueSink_io_deq_bits_opcode;
  assign _T_115_bits_param = AsyncQueueSink_io_deq_bits_param;
  assign _T_115_bits_size = AsyncQueueSink_io_deq_bits_size;
  assign _T_115_bits_source = AsyncQueueSink_io_deq_bits_source;
  assign _T_115_bits_sink = AsyncQueueSink_io_deq_bits_sink;
  assign _T_115_bits_data = AsyncQueueSink_io_deq_bits_data;
  assign _T_115_bits_error = AsyncQueueSink_io_deq_bits_error;
endmodule
module AsyncQueueSource_1(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input        io_enq_bits_resumereq,
  input  [9:0] io_enq_bits_hartsel,
  input        io_ridx,
  output       io_widx,
  output       io_mem_0_resumereq,
  output [9:0] io_mem_0_hartsel,
  input        io_sink_reset_n,
  input        io_ridx_valid,
  output       io_widx_valid
);
  wire  sink_ready;
  reg  mem_0_resumereq;
  reg [31:0] _RAND_0;
  reg [9:0] mem_0_hartsel;
  reg [31:0] _RAND_1;
  wire  _T_26;
  wire  _T_28;
  wire  widx_bin_clock;
  wire  widx_bin_reset;
  wire  widx_bin_io_d;
  wire  widx_bin_io_q;
  wire  widx_bin_io_en;
  wire [1:0] _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_37;
  wire  widx;
  wire  ridx_gray_sync_0_clock;
  wire  ridx_gray_sync_0_reset;
  wire  ridx_gray_sync_0_io_d;
  wire  ridx_gray_sync_0_io_q;
  wire  ridx_gray_sync_0_io_en;
  wire  ridx_gray_sync_1_clock;
  wire  ridx_gray_sync_1_reset;
  wire  ridx_gray_sync_1_io_d;
  wire  ridx_gray_sync_1_io_q;
  wire  ridx_gray_sync_1_io_en;
  wire  ridx_gray_sync_2_clock;
  wire  ridx_gray_sync_2_reset;
  wire  ridx_gray_sync_2_io_d;
  wire  ridx_gray_sync_2_io_q;
  wire  ridx_gray_sync_2_io_en;
  wire  _T_42;
  wire  _T_43;
  wire  ready;
  wire  _GEN_0;
  wire [9:0] _GEN_1;
  wire  ready_reg_clock;
  wire  ready_reg_reset;
  wire  ready_reg_io_d;
  wire  ready_reg_io_q;
  wire  ready_reg_io_en;
  wire  ready_reg_1;
  wire  _T_48;
  wire  widx_gray_clock;
  wire  widx_gray_reset;
  wire  widx_gray_io_d;
  wire  widx_gray_io_q;
  wire  widx_gray_io_en;
  wire  AsyncValidSync_clock;
  wire  AsyncValidSync_reset;
  wire  AsyncValidSync_io_in;
  wire  AsyncValidSync_io_out;
  wire  AsyncValidSync_1_clock;
  wire  AsyncValidSync_1_reset;
  wire  AsyncValidSync_1_io_in;
  wire  AsyncValidSync_1_io_out;
  wire  AsyncValidSync_2_clock;
  wire  AsyncValidSync_2_reset;
  wire  AsyncValidSync_2_io_in;
  wire  AsyncValidSync_2_io_out;
  wire  _T_52;
  wire  _T_53;
  AsyncResetRegVec_1 widx_bin (
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_0 (
    .clock(ridx_gray_sync_0_clock),
    .reset(ridx_gray_sync_0_reset),
    .io_d(ridx_gray_sync_0_io_d),
    .io_q(ridx_gray_sync_0_io_q),
    .io_en(ridx_gray_sync_0_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_1 (
    .clock(ridx_gray_sync_1_clock),
    .reset(ridx_gray_sync_1_reset),
    .io_d(ridx_gray_sync_1_io_d),
    .io_q(ridx_gray_sync_1_io_q),
    .io_en(ridx_gray_sync_1_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_2 (
    .clock(ridx_gray_sync_2_clock),
    .reset(ridx_gray_sync_2_reset),
    .io_d(ridx_gray_sync_2_io_d),
    .io_q(ridx_gray_sync_2_io_q),
    .io_en(ridx_gray_sync_2_io_en)
  );
  AsyncResetRegVec_1 ready_reg (
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_1 widx_gray (
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync (
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 (
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 (
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign io_enq_ready = _T_48;
  assign io_widx = widx_gray_io_q;
  assign io_mem_0_resumereq = mem_0_resumereq;
  assign io_mem_0_hartsel = mem_0_hartsel;
  assign io_widx_valid = AsyncValidSync_io_out;
  assign sink_ready = AsyncValidSync_2_io_out;
  assign _T_26 = io_enq_ready & io_enq_valid;
  assign _T_28 = sink_ready == 1'h0;
  assign widx_bin_clock = clock;
  assign widx_bin_reset = reset;
  assign widx_bin_io_d = _T_35;
  assign widx_bin_io_en = 1'h1;
  assign _T_33 = widx_bin_io_q + _T_26;
  assign _T_34 = _T_33[0:0];
  assign _T_35 = _T_28 ? 1'h0 : _T_34;
  assign _T_37 = _T_35 >> 1'h1;
  assign widx = _T_35 ^ _T_37;
  assign ridx_gray_sync_0_clock = clock;
  assign ridx_gray_sync_0_reset = reset;
  assign ridx_gray_sync_0_io_d = ridx_gray_sync_1_io_q;
  assign ridx_gray_sync_0_io_en = 1'h1;
  assign ridx_gray_sync_1_clock = clock;
  assign ridx_gray_sync_1_reset = reset;
  assign ridx_gray_sync_1_io_d = ridx_gray_sync_2_io_q;
  assign ridx_gray_sync_1_io_en = 1'h1;
  assign ridx_gray_sync_2_clock = clock;
  assign ridx_gray_sync_2_reset = reset;
  assign ridx_gray_sync_2_io_d = io_ridx;
  assign ridx_gray_sync_2_io_en = 1'h1;
  assign _T_42 = ridx_gray_sync_0_io_q ^ 1'h1;
  assign _T_43 = widx != _T_42;
  assign ready = sink_ready & _T_43;
  assign _GEN_0 = _T_26 ? io_enq_bits_resumereq : mem_0_resumereq;
  assign _GEN_1 = _T_26 ? io_enq_bits_hartsel : mem_0_hartsel;
  assign ready_reg_clock = clock;
  assign ready_reg_reset = reset;
  assign ready_reg_io_d = ready;
  assign ready_reg_io_en = 1'h1;
  assign ready_reg_1 = ready_reg_io_q;
  assign _T_48 = ready_reg_1 & sink_ready;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = widx;
  assign widx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_53;
  assign AsyncValidSync_io_in = 1'h1;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_53;
  assign AsyncValidSync_1_io_in = io_ridx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign _T_52 = io_sink_reset_n == 1'h0;
  assign _T_53 = reset | _T_52;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  mem_0_resumereq = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0_hartsel = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_26) begin
      mem_0_resumereq <= io_enq_bits_resumereq;
    end
    if (_T_26) begin
      mem_0_hartsel <= io_enq_bits_hartsel;
    end
  end
endmodule
module TLDebugModuleOuterAsync_dmOuter(
  input         clock,
  input         reset,
  output        io_debugInterrupts_0_0,
  output [2:0]  io_dmiInner_0_a_mem_0_opcode,
  output [1:0]  io_dmiInner_0_a_mem_0_size,
  output        io_dmiInner_0_a_mem_0_source,
  output [8:0]  io_dmiInner_0_a_mem_0_address,
  output [3:0]  io_dmiInner_0_a_mem_0_mask,
  output [31:0] io_dmiInner_0_a_mem_0_data,
  input         io_dmiInner_0_a_ridx,
  output        io_dmiInner_0_a_widx,
  input         io_dmiInner_0_a_ridx_valid,
  output        io_dmiInner_0_a_widx_valid,
  output        io_dmiInner_0_a_source_reset_n,
  input         io_dmiInner_0_a_sink_reset_n,
  input  [2:0]  io_dmiInner_0_d_mem_0_opcode,
  input  [1:0]  io_dmiInner_0_d_mem_0_param,
  input  [1:0]  io_dmiInner_0_d_mem_0_size,
  input         io_dmiInner_0_d_mem_0_source,
  input         io_dmiInner_0_d_mem_0_sink,
  input  [31:0] io_dmiInner_0_d_mem_0_data,
  input         io_dmiInner_0_d_mem_0_error,
  output        io_dmiInner_0_d_ridx,
  input         io_dmiInner_0_d_widx,
  output        io_dmiInner_0_d_ridx_valid,
  input         io_dmiInner_0_d_widx_valid,
  input         io_dmiInner_0_d_source_reset_n,
  output        io_dmiInner_0_d_sink_reset_n,
  output        io_dmi_req_ready,
  input         io_dmi_req_valid,
  input  [6:0]  io_dmi_req_bits_addr,
  input  [31:0] io_dmi_req_bits_data,
  input  [1:0]  io_dmi_req_bits_op,
  input         io_dmi_resp_ready,
  output        io_dmi_resp_valid,
  output [31:0] io_dmi_resp_bits_data,
  output [1:0]  io_dmi_resp_bits_resp,
  output        io_ctrl_ndreset,
  output        io_ctrl_dmactive,
  output        io_innerCtrl_mem_0_resumereq,
  output [9:0]  io_innerCtrl_mem_0_hartsel,
  input         io_innerCtrl_ridx,
  output        io_innerCtrl_widx,
  input         io_innerCtrl_ridx_valid,
  output        io_innerCtrl_widx_valid,
  output        io_innerCtrl_source_reset_n,
  input         io_innerCtrl_sink_reset_n
);
  wire  dmi2tl_io_dmi_req_ready;
  wire  dmi2tl_io_dmi_req_valid;
  wire [6:0] dmi2tl_io_dmi_req_bits_addr;
  wire [31:0] dmi2tl_io_dmi_req_bits_data;
  wire [1:0] dmi2tl_io_dmi_req_bits_op;
  wire  dmi2tl_io_dmi_resp_ready;
  wire  dmi2tl_io_dmi_resp_valid;
  wire [31:0] dmi2tl_io_dmi_resp_bits_data;
  wire [1:0] dmi2tl_io_dmi_resp_bits_resp;
  wire  dmi2tl_io_out_0_a_ready;
  wire  dmi2tl_io_out_0_a_valid;
  wire [2:0] dmi2tl_io_out_0_a_bits_opcode;
  wire [1:0] dmi2tl_io_out_0_a_bits_size;
  wire  dmi2tl_io_out_0_a_bits_source;
  wire [8:0] dmi2tl_io_out_0_a_bits_address;
  wire [3:0] dmi2tl_io_out_0_a_bits_mask;
  wire [31:0] dmi2tl_io_out_0_a_bits_data;
  wire  dmi2tl_io_out_0_d_ready;
  wire  dmi2tl_io_out_0_d_valid;
  wire [31:0] dmi2tl_io_out_0_d_bits_data;
  wire  dmi2tl_io_out_0_d_bits_error;
  wire  dmiXbar_clock;
  wire  dmiXbar_reset;
  wire  dmiXbar_io_in_0_a_ready;
  wire  dmiXbar_io_in_0_a_valid;
  wire [2:0] dmiXbar_io_in_0_a_bits_opcode;
  wire [1:0] dmiXbar_io_in_0_a_bits_size;
  wire  dmiXbar_io_in_0_a_bits_source;
  wire [8:0] dmiXbar_io_in_0_a_bits_address;
  wire [3:0] dmiXbar_io_in_0_a_bits_mask;
  wire [31:0] dmiXbar_io_in_0_a_bits_data;
  wire  dmiXbar_io_in_0_d_ready;
  wire  dmiXbar_io_in_0_d_valid;
  wire [31:0] dmiXbar_io_in_0_d_bits_data;
  wire  dmiXbar_io_in_0_d_bits_error;
  wire  dmiXbar_io_out_1_a_ready;
  wire  dmiXbar_io_out_1_a_valid;
  wire [2:0] dmiXbar_io_out_1_a_bits_opcode;
  wire [1:0] dmiXbar_io_out_1_a_bits_size;
  wire  dmiXbar_io_out_1_a_bits_source;
  wire [8:0] dmiXbar_io_out_1_a_bits_address;
  wire [3:0] dmiXbar_io_out_1_a_bits_mask;
  wire [31:0] dmiXbar_io_out_1_a_bits_data;
  wire  dmiXbar_io_out_1_d_ready;
  wire  dmiXbar_io_out_1_d_valid;
  wire [2:0] dmiXbar_io_out_1_d_bits_opcode;
  wire [1:0] dmiXbar_io_out_1_d_bits_param;
  wire [1:0] dmiXbar_io_out_1_d_bits_size;
  wire  dmiXbar_io_out_1_d_bits_source;
  wire  dmiXbar_io_out_1_d_bits_sink;
  wire [31:0] dmiXbar_io_out_1_d_bits_data;
  wire  dmiXbar_io_out_1_d_bits_error;
  wire  dmiXbar_io_out_0_a_ready;
  wire  dmiXbar_io_out_0_a_valid;
  wire [2:0] dmiXbar_io_out_0_a_bits_opcode;
  wire [1:0] dmiXbar_io_out_0_a_bits_size;
  wire  dmiXbar_io_out_0_a_bits_source;
  wire [6:0] dmiXbar_io_out_0_a_bits_address;
  wire [3:0] dmiXbar_io_out_0_a_bits_mask;
  wire [31:0] dmiXbar_io_out_0_a_bits_data;
  wire  dmiXbar_io_out_0_d_ready;
  wire  dmiXbar_io_out_0_d_valid;
  wire [2:0] dmiXbar_io_out_0_d_bits_opcode;
  wire [1:0] dmiXbar_io_out_0_d_bits_param;
  wire [1:0] dmiXbar_io_out_0_d_bits_size;
  wire  dmiXbar_io_out_0_d_bits_source;
  wire  dmiXbar_io_out_0_d_bits_sink;
  wire [31:0] dmiXbar_io_out_0_d_bits_data;
  wire  dmiXbar_io_out_0_d_bits_error;
  wire  dmOuter_clock;
  wire  dmOuter_reset;
  wire  dmOuter_io_debugInterrupts_0_0;
  wire  dmOuter_io_ctrl_ndreset;
  wire  dmOuter_io_ctrl_dmactive;
  wire  dmOuter_io_tlIn_0_a_ready;
  wire  dmOuter_io_tlIn_0_a_valid;
  wire [2:0] dmOuter_io_tlIn_0_a_bits_opcode;
  wire [1:0] dmOuter_io_tlIn_0_a_bits_size;
  wire  dmOuter_io_tlIn_0_a_bits_source;
  wire [6:0] dmOuter_io_tlIn_0_a_bits_address;
  wire [3:0] dmOuter_io_tlIn_0_a_bits_mask;
  wire [31:0] dmOuter_io_tlIn_0_a_bits_data;
  wire  dmOuter_io_tlIn_0_d_ready;
  wire  dmOuter_io_tlIn_0_d_valid;
  wire [2:0] dmOuter_io_tlIn_0_d_bits_opcode;
  wire [1:0] dmOuter_io_tlIn_0_d_bits_param;
  wire [1:0] dmOuter_io_tlIn_0_d_bits_size;
  wire  dmOuter_io_tlIn_0_d_bits_source;
  wire  dmOuter_io_tlIn_0_d_bits_sink;
  wire [31:0] dmOuter_io_tlIn_0_d_bits_data;
  wire  dmOuter_io_tlIn_0_d_bits_error;
  wire  dmOuter_io_innerCtrl_valid;
  wire  dmOuter_io_innerCtrl_bits_resumereq;
  wire [9:0] dmOuter_io_innerCtrl_bits_hartsel;
  wire  dmInner_TLAsyncCrossingSource_clock;
  wire  dmInner_TLAsyncCrossingSource_reset;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_a_ready;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_a_valid;
  wire [2:0] dmInner_TLAsyncCrossingSource_io_in_0_a_bits_opcode;
  wire [1:0] dmInner_TLAsyncCrossingSource_io_in_0_a_bits_size;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_a_bits_source;
  wire [8:0] dmInner_TLAsyncCrossingSource_io_in_0_a_bits_address;
  wire [3:0] dmInner_TLAsyncCrossingSource_io_in_0_a_bits_mask;
  wire [31:0] dmInner_TLAsyncCrossingSource_io_in_0_a_bits_data;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_d_ready;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_d_valid;
  wire [2:0] dmInner_TLAsyncCrossingSource_io_in_0_d_bits_opcode;
  wire [1:0] dmInner_TLAsyncCrossingSource_io_in_0_d_bits_param;
  wire [1:0] dmInner_TLAsyncCrossingSource_io_in_0_d_bits_size;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_d_bits_source;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_d_bits_sink;
  wire [31:0] dmInner_TLAsyncCrossingSource_io_in_0_d_bits_data;
  wire  dmInner_TLAsyncCrossingSource_io_in_0_d_bits_error;
  wire [2:0] dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_opcode;
  wire [1:0] dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_size;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_source;
  wire [8:0] dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_address;
  wire [3:0] dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_mask;
  wire [31:0] dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_data;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_ridx;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_widx;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_ridx_valid;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_widx_valid;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_source_reset_n;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_a_sink_reset_n;
  wire [2:0] dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_opcode;
  wire [1:0] dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_param;
  wire [1:0] dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_size;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_source;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_sink;
  wire [31:0] dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_data;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_error;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_ridx;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_widx;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_ridx_valid;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_widx_valid;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_source_reset_n;
  wire  dmInner_TLAsyncCrossingSource_io_out_0_d_sink_reset_n;
  wire  AsyncQueueSource_clock;
  wire  AsyncQueueSource_reset;
  wire  AsyncQueueSource_io_enq_ready;
  wire  AsyncQueueSource_io_enq_valid;
  wire  AsyncQueueSource_io_enq_bits_resumereq;
  wire [9:0] AsyncQueueSource_io_enq_bits_hartsel;
  wire  AsyncQueueSource_io_ridx;
  wire  AsyncQueueSource_io_widx;
  wire  AsyncQueueSource_io_mem_0_resumereq;
  wire [9:0] AsyncQueueSource_io_mem_0_hartsel;
  wire  AsyncQueueSource_io_sink_reset_n;
  wire  AsyncQueueSource_io_ridx_valid;
  wire  AsyncQueueSource_io_widx_valid;
  wire  _T_86_mem_0_resumereq;
  wire [9:0] _T_86_mem_0_hartsel;
  wire  _T_86_widx;
  wire  _T_86_widx_valid;
  wire  _T_92;
  DMIToTL_dmi2tl dmi2tl (
    .io_dmi_req_ready(dmi2tl_io_dmi_req_ready),
    .io_dmi_req_valid(dmi2tl_io_dmi_req_valid),
    .io_dmi_req_bits_addr(dmi2tl_io_dmi_req_bits_addr),
    .io_dmi_req_bits_data(dmi2tl_io_dmi_req_bits_data),
    .io_dmi_req_bits_op(dmi2tl_io_dmi_req_bits_op),
    .io_dmi_resp_ready(dmi2tl_io_dmi_resp_ready),
    .io_dmi_resp_valid(dmi2tl_io_dmi_resp_valid),
    .io_dmi_resp_bits_data(dmi2tl_io_dmi_resp_bits_data),
    .io_dmi_resp_bits_resp(dmi2tl_io_dmi_resp_bits_resp),
    .io_out_0_a_ready(dmi2tl_io_out_0_a_ready),
    .io_out_0_a_valid(dmi2tl_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(dmi2tl_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(dmi2tl_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(dmi2tl_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(dmi2tl_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(dmi2tl_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(dmi2tl_io_out_0_a_bits_data),
    .io_out_0_d_ready(dmi2tl_io_out_0_d_ready),
    .io_out_0_d_valid(dmi2tl_io_out_0_d_valid),
    .io_out_0_d_bits_data(dmi2tl_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(dmi2tl_io_out_0_d_bits_error)
  );
  TLXbar_dmiXbar dmiXbar (
    .clock(dmiXbar_clock),
    .reset(dmiXbar_reset),
    .io_in_0_a_ready(dmiXbar_io_in_0_a_ready),
    .io_in_0_a_valid(dmiXbar_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(dmiXbar_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(dmiXbar_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(dmiXbar_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(dmiXbar_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(dmiXbar_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(dmiXbar_io_in_0_a_bits_data),
    .io_in_0_d_ready(dmiXbar_io_in_0_d_ready),
    .io_in_0_d_valid(dmiXbar_io_in_0_d_valid),
    .io_in_0_d_bits_data(dmiXbar_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(dmiXbar_io_in_0_d_bits_error),
    .io_out_1_a_ready(dmiXbar_io_out_1_a_ready),
    .io_out_1_a_valid(dmiXbar_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(dmiXbar_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(dmiXbar_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(dmiXbar_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(dmiXbar_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(dmiXbar_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(dmiXbar_io_out_1_a_bits_data),
    .io_out_1_d_ready(dmiXbar_io_out_1_d_ready),
    .io_out_1_d_valid(dmiXbar_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(dmiXbar_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(dmiXbar_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(dmiXbar_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(dmiXbar_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(dmiXbar_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(dmiXbar_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(dmiXbar_io_out_1_d_bits_error),
    .io_out_0_a_ready(dmiXbar_io_out_0_a_ready),
    .io_out_0_a_valid(dmiXbar_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(dmiXbar_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(dmiXbar_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(dmiXbar_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(dmiXbar_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(dmiXbar_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(dmiXbar_io_out_0_a_bits_data),
    .io_out_0_d_ready(dmiXbar_io_out_0_d_ready),
    .io_out_0_d_valid(dmiXbar_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(dmiXbar_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(dmiXbar_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(dmiXbar_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(dmiXbar_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(dmiXbar_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(dmiXbar_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(dmiXbar_io_out_0_d_bits_error)
  );
  TLDebugModuleOuter_dmOuter dmOuter (
    .clock(dmOuter_clock),
    .reset(dmOuter_reset),
    .io_debugInterrupts_0_0(dmOuter_io_debugInterrupts_0_0),
    .io_ctrl_ndreset(dmOuter_io_ctrl_ndreset),
    .io_ctrl_dmactive(dmOuter_io_ctrl_dmactive),
    .io_tlIn_0_a_ready(dmOuter_io_tlIn_0_a_ready),
    .io_tlIn_0_a_valid(dmOuter_io_tlIn_0_a_valid),
    .io_tlIn_0_a_bits_opcode(dmOuter_io_tlIn_0_a_bits_opcode),
    .io_tlIn_0_a_bits_size(dmOuter_io_tlIn_0_a_bits_size),
    .io_tlIn_0_a_bits_source(dmOuter_io_tlIn_0_a_bits_source),
    .io_tlIn_0_a_bits_address(dmOuter_io_tlIn_0_a_bits_address),
    .io_tlIn_0_a_bits_mask(dmOuter_io_tlIn_0_a_bits_mask),
    .io_tlIn_0_a_bits_data(dmOuter_io_tlIn_0_a_bits_data),
    .io_tlIn_0_d_ready(dmOuter_io_tlIn_0_d_ready),
    .io_tlIn_0_d_valid(dmOuter_io_tlIn_0_d_valid),
    .io_tlIn_0_d_bits_opcode(dmOuter_io_tlIn_0_d_bits_opcode),
    .io_tlIn_0_d_bits_param(dmOuter_io_tlIn_0_d_bits_param),
    .io_tlIn_0_d_bits_size(dmOuter_io_tlIn_0_d_bits_size),
    .io_tlIn_0_d_bits_source(dmOuter_io_tlIn_0_d_bits_source),
    .io_tlIn_0_d_bits_sink(dmOuter_io_tlIn_0_d_bits_sink),
    .io_tlIn_0_d_bits_data(dmOuter_io_tlIn_0_d_bits_data),
    .io_tlIn_0_d_bits_error(dmOuter_io_tlIn_0_d_bits_error),
    .io_innerCtrl_valid(dmOuter_io_innerCtrl_valid),
    .io_innerCtrl_bits_resumereq(dmOuter_io_innerCtrl_bits_resumereq),
    .io_innerCtrl_bits_hartsel(dmOuter_io_innerCtrl_bits_hartsel)
  );
  TLAsyncCrossingSource_dmInner dmInner_TLAsyncCrossingSource (
    .clock(dmInner_TLAsyncCrossingSource_clock),
    .reset(dmInner_TLAsyncCrossingSource_reset),
    .io_in_0_a_ready(dmInner_TLAsyncCrossingSource_io_in_0_a_ready),
    .io_in_0_a_valid(dmInner_TLAsyncCrossingSource_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(dmInner_TLAsyncCrossingSource_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(dmInner_TLAsyncCrossingSource_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(dmInner_TLAsyncCrossingSource_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(dmInner_TLAsyncCrossingSource_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(dmInner_TLAsyncCrossingSource_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(dmInner_TLAsyncCrossingSource_io_in_0_a_bits_data),
    .io_in_0_d_ready(dmInner_TLAsyncCrossingSource_io_in_0_d_ready),
    .io_in_0_d_valid(dmInner_TLAsyncCrossingSource_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(dmInner_TLAsyncCrossingSource_io_in_0_d_bits_error),
    .io_out_0_a_mem_0_opcode(dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_opcode),
    .io_out_0_a_mem_0_size(dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_size),
    .io_out_0_a_mem_0_source(dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_source),
    .io_out_0_a_mem_0_address(dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_address),
    .io_out_0_a_mem_0_mask(dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_mask),
    .io_out_0_a_mem_0_data(dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_data),
    .io_out_0_a_ridx(dmInner_TLAsyncCrossingSource_io_out_0_a_ridx),
    .io_out_0_a_widx(dmInner_TLAsyncCrossingSource_io_out_0_a_widx),
    .io_out_0_a_ridx_valid(dmInner_TLAsyncCrossingSource_io_out_0_a_ridx_valid),
    .io_out_0_a_widx_valid(dmInner_TLAsyncCrossingSource_io_out_0_a_widx_valid),
    .io_out_0_a_source_reset_n(dmInner_TLAsyncCrossingSource_io_out_0_a_source_reset_n),
    .io_out_0_a_sink_reset_n(dmInner_TLAsyncCrossingSource_io_out_0_a_sink_reset_n),
    .io_out_0_d_mem_0_opcode(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_opcode),
    .io_out_0_d_mem_0_param(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_param),
    .io_out_0_d_mem_0_size(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_size),
    .io_out_0_d_mem_0_source(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_source),
    .io_out_0_d_mem_0_sink(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_sink),
    .io_out_0_d_mem_0_data(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_data),
    .io_out_0_d_mem_0_error(dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_error),
    .io_out_0_d_ridx(dmInner_TLAsyncCrossingSource_io_out_0_d_ridx),
    .io_out_0_d_widx(dmInner_TLAsyncCrossingSource_io_out_0_d_widx),
    .io_out_0_d_ridx_valid(dmInner_TLAsyncCrossingSource_io_out_0_d_ridx_valid),
    .io_out_0_d_widx_valid(dmInner_TLAsyncCrossingSource_io_out_0_d_widx_valid),
    .io_out_0_d_source_reset_n(dmInner_TLAsyncCrossingSource_io_out_0_d_source_reset_n),
    .io_out_0_d_sink_reset_n(dmInner_TLAsyncCrossingSource_io_out_0_d_sink_reset_n)
  );
  AsyncQueueSource_1 AsyncQueueSource (
    .clock(AsyncQueueSource_clock),
    .reset(AsyncQueueSource_reset),
    .io_enq_ready(AsyncQueueSource_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_io_enq_valid),
    .io_enq_bits_resumereq(AsyncQueueSource_io_enq_bits_resumereq),
    .io_enq_bits_hartsel(AsyncQueueSource_io_enq_bits_hartsel),
    .io_ridx(AsyncQueueSource_io_ridx),
    .io_widx(AsyncQueueSource_io_widx),
    .io_mem_0_resumereq(AsyncQueueSource_io_mem_0_resumereq),
    .io_mem_0_hartsel(AsyncQueueSource_io_mem_0_hartsel),
    .io_sink_reset_n(AsyncQueueSource_io_sink_reset_n),
    .io_ridx_valid(AsyncQueueSource_io_ridx_valid),
    .io_widx_valid(AsyncQueueSource_io_widx_valid)
  );
  assign io_debugInterrupts_0_0 = dmOuter_io_debugInterrupts_0_0;
  assign io_dmiInner_0_a_mem_0_opcode = dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_opcode;
  assign io_dmiInner_0_a_mem_0_size = dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_size;
  assign io_dmiInner_0_a_mem_0_source = dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_source;
  assign io_dmiInner_0_a_mem_0_address = dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_address;
  assign io_dmiInner_0_a_mem_0_mask = dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_mask;
  assign io_dmiInner_0_a_mem_0_data = dmInner_TLAsyncCrossingSource_io_out_0_a_mem_0_data;
  assign io_dmiInner_0_a_widx = dmInner_TLAsyncCrossingSource_io_out_0_a_widx;
  assign io_dmiInner_0_a_widx_valid = dmInner_TLAsyncCrossingSource_io_out_0_a_widx_valid;
  assign io_dmiInner_0_a_source_reset_n = dmInner_TLAsyncCrossingSource_io_out_0_a_source_reset_n;
  assign io_dmiInner_0_d_ridx = dmInner_TLAsyncCrossingSource_io_out_0_d_ridx;
  assign io_dmiInner_0_d_ridx_valid = dmInner_TLAsyncCrossingSource_io_out_0_d_ridx_valid;
  assign io_dmiInner_0_d_sink_reset_n = dmInner_TLAsyncCrossingSource_io_out_0_d_sink_reset_n;
  assign io_dmi_req_ready = dmi2tl_io_dmi_req_ready;
  assign io_dmi_resp_valid = dmi2tl_io_dmi_resp_valid;
  assign io_dmi_resp_bits_data = dmi2tl_io_dmi_resp_bits_data;
  assign io_dmi_resp_bits_resp = dmi2tl_io_dmi_resp_bits_resp;
  assign io_ctrl_ndreset = dmOuter_io_ctrl_ndreset;
  assign io_ctrl_dmactive = dmOuter_io_ctrl_dmactive;
  assign io_innerCtrl_mem_0_resumereq = _T_86_mem_0_resumereq;
  assign io_innerCtrl_mem_0_hartsel = _T_86_mem_0_hartsel;
  assign io_innerCtrl_widx = _T_86_widx;
  assign io_innerCtrl_widx_valid = _T_86_widx_valid;
  assign io_innerCtrl_source_reset_n = _T_92;
  assign dmi2tl_io_dmi_req_valid = io_dmi_req_valid;
  assign dmi2tl_io_dmi_req_bits_addr = io_dmi_req_bits_addr;
  assign dmi2tl_io_dmi_req_bits_data = io_dmi_req_bits_data;
  assign dmi2tl_io_dmi_req_bits_op = io_dmi_req_bits_op;
  assign dmi2tl_io_dmi_resp_ready = io_dmi_resp_ready;
  assign dmi2tl_io_out_0_a_ready = dmiXbar_io_in_0_a_ready;
  assign dmi2tl_io_out_0_d_valid = dmiXbar_io_in_0_d_valid;
  assign dmi2tl_io_out_0_d_bits_data = dmiXbar_io_in_0_d_bits_data;
  assign dmi2tl_io_out_0_d_bits_error = dmiXbar_io_in_0_d_bits_error;
  assign dmiXbar_clock = clock;
  assign dmiXbar_reset = reset;
  assign dmiXbar_io_in_0_a_valid = dmi2tl_io_out_0_a_valid;
  assign dmiXbar_io_in_0_a_bits_opcode = dmi2tl_io_out_0_a_bits_opcode;
  assign dmiXbar_io_in_0_a_bits_size = dmi2tl_io_out_0_a_bits_size;
  assign dmiXbar_io_in_0_a_bits_source = dmi2tl_io_out_0_a_bits_source;
  assign dmiXbar_io_in_0_a_bits_address = dmi2tl_io_out_0_a_bits_address;
  assign dmiXbar_io_in_0_a_bits_mask = dmi2tl_io_out_0_a_bits_mask;
  assign dmiXbar_io_in_0_a_bits_data = dmi2tl_io_out_0_a_bits_data;
  assign dmiXbar_io_in_0_d_ready = dmi2tl_io_out_0_d_ready;
  assign dmiXbar_io_out_1_a_ready = dmInner_TLAsyncCrossingSource_io_in_0_a_ready;
  assign dmiXbar_io_out_1_d_valid = dmInner_TLAsyncCrossingSource_io_in_0_d_valid;
  assign dmiXbar_io_out_1_d_bits_opcode = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_opcode;
  assign dmiXbar_io_out_1_d_bits_param = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_param;
  assign dmiXbar_io_out_1_d_bits_size = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_size;
  assign dmiXbar_io_out_1_d_bits_source = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_source;
  assign dmiXbar_io_out_1_d_bits_sink = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_sink;
  assign dmiXbar_io_out_1_d_bits_data = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_data;
  assign dmiXbar_io_out_1_d_bits_error = dmInner_TLAsyncCrossingSource_io_in_0_d_bits_error;
  assign dmiXbar_io_out_0_a_ready = dmOuter_io_tlIn_0_a_ready;
  assign dmiXbar_io_out_0_d_valid = dmOuter_io_tlIn_0_d_valid;
  assign dmiXbar_io_out_0_d_bits_opcode = dmOuter_io_tlIn_0_d_bits_opcode;
  assign dmiXbar_io_out_0_d_bits_param = dmOuter_io_tlIn_0_d_bits_param;
  assign dmiXbar_io_out_0_d_bits_size = dmOuter_io_tlIn_0_d_bits_size;
  assign dmiXbar_io_out_0_d_bits_source = dmOuter_io_tlIn_0_d_bits_source;
  assign dmiXbar_io_out_0_d_bits_sink = dmOuter_io_tlIn_0_d_bits_sink;
  assign dmiXbar_io_out_0_d_bits_data = dmOuter_io_tlIn_0_d_bits_data;
  assign dmiXbar_io_out_0_d_bits_error = dmOuter_io_tlIn_0_d_bits_error;
  assign dmOuter_clock = clock;
  assign dmOuter_reset = reset;
  assign dmOuter_io_tlIn_0_a_valid = dmiXbar_io_out_0_a_valid;
  assign dmOuter_io_tlIn_0_a_bits_opcode = dmiXbar_io_out_0_a_bits_opcode;
  assign dmOuter_io_tlIn_0_a_bits_size = dmiXbar_io_out_0_a_bits_size;
  assign dmOuter_io_tlIn_0_a_bits_source = dmiXbar_io_out_0_a_bits_source;
  assign dmOuter_io_tlIn_0_a_bits_address = dmiXbar_io_out_0_a_bits_address;
  assign dmOuter_io_tlIn_0_a_bits_mask = dmiXbar_io_out_0_a_bits_mask;
  assign dmOuter_io_tlIn_0_a_bits_data = dmiXbar_io_out_0_a_bits_data;
  assign dmOuter_io_tlIn_0_d_ready = dmiXbar_io_out_0_d_ready;
  assign dmInner_TLAsyncCrossingSource_clock = clock;
  assign dmInner_TLAsyncCrossingSource_reset = reset;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_valid = dmiXbar_io_out_1_a_valid;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_bits_opcode = dmiXbar_io_out_1_a_bits_opcode;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_bits_size = dmiXbar_io_out_1_a_bits_size;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_bits_source = dmiXbar_io_out_1_a_bits_source;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_bits_address = dmiXbar_io_out_1_a_bits_address;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_bits_mask = dmiXbar_io_out_1_a_bits_mask;
  assign dmInner_TLAsyncCrossingSource_io_in_0_a_bits_data = dmiXbar_io_out_1_a_bits_data;
  assign dmInner_TLAsyncCrossingSource_io_in_0_d_ready = dmiXbar_io_out_1_d_ready;
  assign dmInner_TLAsyncCrossingSource_io_out_0_a_ridx = io_dmiInner_0_a_ridx;
  assign dmInner_TLAsyncCrossingSource_io_out_0_a_ridx_valid = io_dmiInner_0_a_ridx_valid;
  assign dmInner_TLAsyncCrossingSource_io_out_0_a_sink_reset_n = io_dmiInner_0_a_sink_reset_n;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_opcode = io_dmiInner_0_d_mem_0_opcode;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_param = io_dmiInner_0_d_mem_0_param;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_size = io_dmiInner_0_d_mem_0_size;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_source = io_dmiInner_0_d_mem_0_source;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_sink = io_dmiInner_0_d_mem_0_sink;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_data = io_dmiInner_0_d_mem_0_data;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_mem_0_error = io_dmiInner_0_d_mem_0_error;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_widx = io_dmiInner_0_d_widx;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_widx_valid = io_dmiInner_0_d_widx_valid;
  assign dmInner_TLAsyncCrossingSource_io_out_0_d_source_reset_n = io_dmiInner_0_d_source_reset_n;
  assign AsyncQueueSource_clock = clock;
  assign AsyncQueueSource_reset = reset;
  assign AsyncQueueSource_io_enq_valid = dmOuter_io_innerCtrl_valid;
  assign AsyncQueueSource_io_enq_bits_resumereq = dmOuter_io_innerCtrl_bits_resumereq;
  assign AsyncQueueSource_io_enq_bits_hartsel = dmOuter_io_innerCtrl_bits_hartsel;
  assign AsyncQueueSource_io_ridx = io_innerCtrl_ridx;
  assign AsyncQueueSource_io_sink_reset_n = io_innerCtrl_sink_reset_n;
  assign AsyncQueueSource_io_ridx_valid = io_innerCtrl_ridx_valid;
  assign _T_86_mem_0_resumereq = AsyncQueueSource_io_mem_0_resumereq;
  assign _T_86_mem_0_hartsel = AsyncQueueSource_io_mem_0_hartsel;
  assign _T_86_widx = AsyncQueueSource_io_widx;
  assign _T_86_widx_valid = AsyncQueueSource_io_widx_valid;
  assign _T_92 = AsyncQueueSource_reset == 1'h0;
endmodule
module TLDebugModuleInner_dmInner(
  input         clock,
  input         reset,
  output        io_hart_in_0_a_ready,
  input         io_hart_in_0_a_valid,
  input  [2:0]  io_hart_in_0_a_bits_opcode,
  input  [1:0]  io_hart_in_0_a_bits_size,
  input  [9:0]  io_hart_in_0_a_bits_source,
  input  [11:0] io_hart_in_0_a_bits_address,
  input  [3:0]  io_hart_in_0_a_bits_mask,
  input  [31:0] io_hart_in_0_a_bits_data,
  input         io_hart_in_0_d_ready,
  output        io_hart_in_0_d_valid,
  output [2:0]  io_hart_in_0_d_bits_opcode,
  output [1:0]  io_hart_in_0_d_bits_param,
  output [1:0]  io_hart_in_0_d_bits_size,
  output [9:0]  io_hart_in_0_d_bits_source,
  output        io_hart_in_0_d_bits_sink,
  output [31:0] io_hart_in_0_d_bits_data,
  output        io_hart_in_0_d_bits_error,
  output        io_dmi_in_0_a_ready,
  input         io_dmi_in_0_a_valid,
  input  [2:0]  io_dmi_in_0_a_bits_opcode,
  input  [1:0]  io_dmi_in_0_a_bits_size,
  input         io_dmi_in_0_a_bits_source,
  input  [8:0]  io_dmi_in_0_a_bits_address,
  input  [3:0]  io_dmi_in_0_a_bits_mask,
  input  [31:0] io_dmi_in_0_a_bits_data,
  input         io_dmi_in_0_d_ready,
  output        io_dmi_in_0_d_valid,
  output [2:0]  io_dmi_in_0_d_bits_opcode,
  output [1:0]  io_dmi_in_0_d_bits_param,
  output [1:0]  io_dmi_in_0_d_bits_size,
  output        io_dmi_in_0_d_bits_source,
  output        io_dmi_in_0_d_bits_sink,
  output [31:0] io_dmi_in_0_d_bits_data,
  output        io_dmi_in_0_d_bits_error,
  input         io_dmactive,
  output        io_innerCtrl_ready,
  input         io_innerCtrl_valid,
  input         io_innerCtrl_bits_resumereq,
  input  [9:0]  io_innerCtrl_bits_hartsel,
  input         io_debugUnavail_0
);
  reg  haltedBitRegs_0;
  reg [31:0] _RAND_0;
  reg  resumeReqRegs_0;
  reg [31:0] _RAND_1;
  reg [9:0] selectedHartReg;
  reg [31:0] _RAND_2;
  wire  _T_1197;
  wire [9:0] _GEN_14;
  wire  _T_1246;
  wire  _T_1254;
  wire  _T_1255;
  wire  _T_1265;
  wire  _T_1266;
  wire  _T_1267;
  wire  _T_1276;
  wire  _T_1277;
  wire  resumereq;
  wire  _T_1285;
  wire  _T_1286;
  wire  _T_1287;
  wire [31:0] haltedStatus_0;
  wire  haltedSummary;
  wire [31:0] _T_1323;
  wire  _T_1324;
  wire  _T_1325;
  wire  _T_1326;
  wire  _T_1327;
  wire  _T_1328;
  wire  _T_1329;
  wire  _T_1330;
  wire  _T_1331;
  wire  _T_1332;
  wire  _T_1333;
  wire  _T_1334;
  wire  _T_1335;
  wire  _T_1336;
  wire  _T_1337;
  wire  _T_1338;
  wire  _T_1339;
  wire  _T_1340;
  wire  _T_1341;
  wire  _T_1342;
  wire  _T_1343;
  wire  _T_1344;
  wire  _T_1345;
  wire  _T_1346;
  wire  _T_1347;
  wire  _T_1348;
  wire  _T_1349;
  wire  _T_1350;
  wire  _T_1351;
  wire  _T_1352;
  wire  _T_1353;
  wire  _T_1354;
  wire  _T_1355;
  reg [2:0] ABSTRACTCSReg_reserved0;
  reg [31:0] _RAND_3;
  reg [4:0] ABSTRACTCSReg_progsize;
  reg [31:0] _RAND_4;
  reg [10:0] ABSTRACTCSReg_reserved1;
  reg [31:0] _RAND_5;
  reg  ABSTRACTCSReg_reserved2;
  reg [31:0] _RAND_6;
  reg [2:0] ABSTRACTCSReg_cmderr;
  reg [31:0] _RAND_7;
  reg [2:0] ABSTRACTCSReg_reserved3;
  reg [31:0] _RAND_8;
  reg [4:0] ABSTRACTCSReg_datacount;
  reg [31:0] _RAND_9;
  wire [2:0] _T_1382;
  wire  ABSTRACTCSWrEn;
  wire  _T_1403;
  wire [2:0] _GEN_23;
  wire [4:0] _GEN_24;
  wire [10:0] _GEN_25;
  wire  _GEN_27;
  wire [2:0] _GEN_28;
  wire [2:0] _GEN_29;
  wire [4:0] _GEN_30;
  wire  _T_1405;
  wire [2:0] _GEN_31;
  wire  _T_1408;
  wire  _T_1409;
  wire [2:0] _GEN_32;
  wire  _T_1414;
  wire  _T_1415;
  wire  _T_1416;
  wire [2:0] _GEN_33;
  wire  _T_1424;
  wire  _T_1425;
  wire  _T_1426;
  wire [2:0] _GEN_34;
  wire  _T_1437;
  wire  _T_1438;
  wire [2:0] _T_1439;
  wire [2:0] _T_1440;
  wire [2:0] _GEN_35;
  wire [2:0] _GEN_36;
  wire [2:0] _GEN_37;
  reg [15:0] ABSTRACTAUTOReg_autoexecprogbuf;
  reg [31:0] _RAND_10;
  reg [3:0] ABSTRACTAUTOReg_reserved0;
  reg [31:0] _RAND_11;
  reg [11:0] ABSTRACTAUTOReg_autoexecdata;
  reg [31:0] _RAND_12;
  wire [11:0] _T_1460;
  wire [15:0] _T_1462;
  wire  ABSTRACTAUTOWrEn;
  wire [15:0] _GEN_38;
  wire [3:0] _GEN_39;
  wire [11:0] _GEN_40;
  wire  _T_1473;
  wire [11:0] _T_1477;
  wire [15:0] _GEN_41;
  wire [11:0] _GEN_42;
  wire  _T_1519;
  wire  _T_1520;
  wire  _T_1521;
  wire  _T_1522;
  wire  _T_1984;
  wire  _T_1985;
  wire  _T_1986;
  wire  _T_1987;
  wire  _T_1988;
  wire  _T_1989;
  wire  _T_1990;
  wire  _T_1991;
  wire  _T_1992;
  wire  _T_1993;
  wire  _T_1994;
  wire  _T_1995;
  wire  _T_1996;
  wire  _T_1997;
  wire  _T_1998;
  wire  _T_1999;
  wire  _T_2000;
  wire  _T_2001;
  wire  _T_2002;
  wire  _T_2003;
  wire  _T_2004;
  wire  _T_2005;
  wire  _T_2006;
  wire  _T_2007;
  wire  _T_2008;
  wire  _T_2009;
  wire  _T_2010;
  wire  _T_2011;
  wire  _T_2012;
  wire  _T_2013;
  wire  _T_2014;
  wire  _T_2015;
  wire  _T_2016;
  wire  _T_2017;
  wire  _T_2018;
  wire  _T_2019;
  wire  _T_2020;
  wire  _T_2021;
  wire  _T_2022;
  wire  _T_2023;
  wire  _T_2024;
  wire  _T_2025;
  wire  _T_2026;
  wire  _T_2027;
  wire  _T_2028;
  wire  _T_2029;
  wire  _T_2030;
  wire  _T_2031;
  wire  _T_2032;
  wire  _T_2033;
  wire  _T_2034;
  wire  _T_2035;
  wire  _T_2036;
  wire  _T_2037;
  wire  _T_2038;
  wire  _T_2039;
  wire  _T_2040;
  wire  _T_2041;
  wire  _T_2042;
  wire  _T_2043;
  wire  _T_2044;
  wire  _T_2045;
  wire  _T_2046;
  wire  _T_2047;
  wire  _T_2048;
  wire  _T_2049;
  wire  dmiAbstractDataAccess;
  wire  _T_2050;
  wire  _T_2051;
  wire  _T_2052;
  wire  _T_2053;
  wire  _T_2054;
  wire  _T_2055;
  wire  _T_2056;
  wire  _T_2057;
  wire  _T_2058;
  wire  _T_2059;
  wire  _T_2060;
  wire  _T_2061;
  wire  _T_2062;
  wire  _T_2063;
  wire  _T_2064;
  wire  _T_2065;
  wire  _T_2066;
  wire  _T_2067;
  wire  _T_2068;
  wire  _T_2069;
  wire  _T_2070;
  wire  _T_2071;
  wire  _T_2072;
  wire  _T_2073;
  wire  _T_2074;
  wire  _T_2075;
  wire  _T_2076;
  wire  _T_2077;
  wire  _T_2078;
  wire  _T_2079;
  wire  _T_2080;
  wire  _T_2081;
  wire  _T_2082;
  wire  _T_2083;
  wire  _T_2084;
  wire  _T_2085;
  wire  _T_2086;
  wire  _T_2087;
  wire  _T_2088;
  wire  _T_2089;
  wire  _T_2090;
  wire  _T_2091;
  wire  _T_2092;
  wire  _T_2093;
  wire  _T_2094;
  wire  _T_2095;
  wire  _T_2096;
  wire  _T_2097;
  wire  _T_2098;
  wire  _T_2099;
  wire  _T_2100;
  wire  _T_2101;
  wire  _T_2102;
  wire  _T_2103;
  wire  _T_2104;
  wire  _T_2105;
  wire  _T_2106;
  wire  _T_2107;
  wire  _T_2108;
  wire  _T_2109;
  wire  _T_2110;
  wire  _T_2111;
  wire  dmiProgramBufferAccess;
  wire  _T_2257;
  wire  _T_2269;
  wire  _T_2270;
  wire  _T_2271;
  wire  _T_2272;
  wire  _T_2273;
  wire  _T_2274;
  wire  _T_2275;
  wire  _T_2276;
  wire  _T_2277;
  wire  _T_2278;
  wire  _T_2279;
  wire  _T_2280;
  wire  _T_2281;
  wire  _T_2282;
  wire  _T_2283;
  wire  _T_2284;
  wire  _T_2285;
  wire  _T_2286;
  wire  _T_2287;
  wire  _T_2288;
  wire  _T_2289;
  wire  _T_2290;
  wire  _T_2291;
  wire  _T_2292;
  wire  _T_2293;
  wire  _T_2294;
  wire  _T_2295;
  wire  _T_2296;
  wire  _T_2297;
  wire  _T_2298;
  wire  _T_2299;
  wire  _T_2300;
  wire  _T_2301;
  wire  _T_2302;
  wire  _T_2303;
  wire  _T_2304;
  wire  _T_2305;
  wire  _T_2306;
  wire  _T_2307;
  wire  _T_2308;
  wire  _T_2309;
  wire  _T_2310;
  wire  _T_2311;
  wire  _T_2312;
  wire  _T_2313;
  wire  _T_2314;
  wire  _T_2315;
  wire  _T_2316;
  wire  autoexec;
  reg [7:0] COMMANDRdData_cmdtype;
  reg [31:0] _RAND_13;
  reg [23:0] COMMANDRdData_control;
  reg [31:0] _RAND_14;
  wire [23:0] _T_2334;
  wire [7:0] _T_2335;
  wire  COMMANDWrEn;
  wire [7:0] _GEN_43;
  wire [23:0] _GEN_44;
  wire [7:0] _GEN_45;
  wire [23:0] _GEN_46;
  wire [7:0] _GEN_47;
  wire [23:0] _GEN_48;
  reg [7:0] abstractDataMem_0;
  reg [31:0] _RAND_15;
  reg [7:0] abstractDataMem_1;
  reg [31:0] _RAND_16;
  reg [7:0] abstractDataMem_2;
  reg [31:0] _RAND_17;
  reg [7:0] abstractDataMem_3;
  reg [31:0] _RAND_18;
  reg [7:0] programBufferMem_0;
  reg [31:0] _RAND_19;
  reg [7:0] programBufferMem_1;
  reg [31:0] _RAND_20;
  reg [7:0] programBufferMem_2;
  reg [31:0] _RAND_21;
  reg [7:0] programBufferMem_3;
  reg [31:0] _RAND_22;
  reg [7:0] programBufferMem_4;
  reg [31:0] _RAND_23;
  reg [7:0] programBufferMem_5;
  reg [31:0] _RAND_24;
  reg [7:0] programBufferMem_6;
  reg [31:0] _RAND_25;
  reg [7:0] programBufferMem_7;
  reg [31:0] _RAND_26;
  reg [7:0] programBufferMem_8;
  reg [31:0] _RAND_27;
  reg [7:0] programBufferMem_9;
  reg [31:0] _RAND_28;
  reg [7:0] programBufferMem_10;
  reg [31:0] _RAND_29;
  reg [7:0] programBufferMem_11;
  reg [31:0] _RAND_30;
  reg [7:0] programBufferMem_12;
  reg [31:0] _RAND_31;
  reg [7:0] programBufferMem_13;
  reg [31:0] _RAND_32;
  reg [7:0] programBufferMem_14;
  reg [31:0] _RAND_33;
  reg [7:0] programBufferMem_15;
  reg [31:0] _RAND_34;
  reg [7:0] programBufferMem_16;
  reg [31:0] _RAND_35;
  reg [7:0] programBufferMem_17;
  reg [31:0] _RAND_36;
  reg [7:0] programBufferMem_18;
  reg [31:0] _RAND_37;
  reg [7:0] programBufferMem_19;
  reg [31:0] _RAND_38;
  reg [7:0] programBufferMem_20;
  reg [31:0] _RAND_39;
  reg [7:0] programBufferMem_21;
  reg [31:0] _RAND_40;
  reg [7:0] programBufferMem_22;
  reg [31:0] _RAND_41;
  reg [7:0] programBufferMem_23;
  reg [31:0] _RAND_42;
  reg [7:0] programBufferMem_24;
  reg [31:0] _RAND_43;
  reg [7:0] programBufferMem_25;
  reg [31:0] _RAND_44;
  reg [7:0] programBufferMem_26;
  reg [31:0] _RAND_45;
  reg [7:0] programBufferMem_27;
  reg [31:0] _RAND_46;
  reg [7:0] programBufferMem_28;
  reg [31:0] _RAND_47;
  reg [7:0] programBufferMem_29;
  reg [31:0] _RAND_48;
  reg [7:0] programBufferMem_30;
  reg [31:0] _RAND_49;
  reg [7:0] programBufferMem_31;
  reg [31:0] _RAND_50;
  reg [7:0] programBufferMem_32;
  reg [31:0] _RAND_51;
  reg [7:0] programBufferMem_33;
  reg [31:0] _RAND_52;
  reg [7:0] programBufferMem_34;
  reg [31:0] _RAND_53;
  reg [7:0] programBufferMem_35;
  reg [31:0] _RAND_54;
  reg [7:0] programBufferMem_36;
  reg [31:0] _RAND_55;
  reg [7:0] programBufferMem_37;
  reg [31:0] _RAND_56;
  reg [7:0] programBufferMem_38;
  reg [31:0] _RAND_57;
  reg [7:0] programBufferMem_39;
  reg [31:0] _RAND_58;
  reg [7:0] programBufferMem_40;
  reg [31:0] _RAND_59;
  reg [7:0] programBufferMem_41;
  reg [31:0] _RAND_60;
  reg [7:0] programBufferMem_42;
  reg [31:0] _RAND_61;
  reg [7:0] programBufferMem_43;
  reg [31:0] _RAND_62;
  reg [7:0] programBufferMem_44;
  reg [31:0] _RAND_63;
  reg [7:0] programBufferMem_45;
  reg [31:0] _RAND_64;
  reg [7:0] programBufferMem_46;
  reg [31:0] _RAND_65;
  reg [7:0] programBufferMem_47;
  reg [31:0] _RAND_66;
  reg [7:0] programBufferMem_48;
  reg [31:0] _RAND_67;
  reg [7:0] programBufferMem_49;
  reg [31:0] _RAND_68;
  reg [7:0] programBufferMem_50;
  reg [31:0] _RAND_69;
  reg [7:0] programBufferMem_51;
  reg [31:0] _RAND_70;
  reg [7:0] programBufferMem_52;
  reg [31:0] _RAND_71;
  reg [7:0] programBufferMem_53;
  reg [31:0] _RAND_72;
  reg [7:0] programBufferMem_54;
  reg [31:0] _RAND_73;
  reg [7:0] programBufferMem_55;
  reg [31:0] _RAND_74;
  reg [7:0] programBufferMem_56;
  reg [31:0] _RAND_75;
  reg [7:0] programBufferMem_57;
  reg [31:0] _RAND_76;
  reg [7:0] programBufferMem_58;
  reg [31:0] _RAND_77;
  reg [7:0] programBufferMem_59;
  reg [31:0] _RAND_78;
  reg [7:0] programBufferMem_60;
  reg [31:0] _RAND_79;
  reg [7:0] programBufferMem_61;
  reg [31:0] _RAND_80;
  reg [7:0] programBufferMem_62;
  reg [31:0] _RAND_81;
  reg [7:0] programBufferMem_63;
  reg [31:0] _RAND_82;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _T_2786;
  wire  _GEN_51;
  wire  _GEN_52;
  wire  _T_2789;
  wire  _T_2790;
  wire  _T_2792;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire [1:0] _T_2806;
  wire [3:0] _T_2807;
  wire [9:0] _T_2808;
  wire [1:0] _T_2809;
  wire [1:0] _T_2810;
  wire [3:0] _T_2811;
  wire [1:0] _T_2812;
  wire [14:0] _T_2813;
  wire [15:0] _T_2814;
  wire [17:0] _T_2815;
  wire [21:0] _T_2816;
  wire [31:0] _T_2817;
  wire [1:0] _T_2823;
  wire [1:0] _T_2824;
  wire [3:0] _T_2825;
  wire [1:0] _T_2826;
  wire [1:0] _T_2827;
  wire [3:0] _T_2828;
  wire [7:0] _T_2829;
  wire [1:0] _T_2830;
  wire [1:0] _T_2831;
  wire [3:0] _T_2832;
  wire [1:0] _T_2833;
  wire [1:0] _T_2834;
  wire [3:0] _T_2835;
  wire [7:0] _T_2836;
  wire [15:0] _T_2837;
  wire [1:0] _T_2838;
  wire [1:0] _T_2839;
  wire [3:0] _T_2840;
  wire [1:0] _T_2841;
  wire [1:0] _T_2842;
  wire [3:0] _T_2843;
  wire [7:0] _T_2844;
  wire [1:0] _T_2845;
  wire [1:0] _T_2846;
  wire [3:0] _T_2847;
  wire [1:0] _T_2848;
  wire [1:0] _T_2849;
  wire [3:0] _T_2850;
  wire [7:0] _T_2851;
  wire [15:0] _T_2852;
  wire [31:0] _T_2853;
  wire [7:0] _T_2854;
  wire [3:0] _T_2855;
  wire [11:0] _T_2856;
  wire [11:0] _T_2857;
  wire [7:0] _T_2858;
  wire [19:0] _T_2859;
  wire [31:0] _T_2860;
  wire [19:0] _T_2861;
  wire [31:0] _T_2862;
  wire [31:0] _T_2863;
  wire  _T_2874;
  wire [6:0] _T_2875;
  wire [2:0] _T_2876;
  wire [6:0] _T_2962;
  wire [6:0] _T_2963;
  wire  _T_2965;
  wire [6:0] _T_2971;
  wire [6:0] _T_2972;
  wire  _T_2974;
  wire [6:0] _T_2980;
  wire [6:0] _T_2981;
  wire  _T_2983;
  wire [6:0] _T_2989;
  wire [6:0] _T_2990;
  wire  _T_2992;
  wire [6:0] _T_2998;
  wire [6:0] _T_2999;
  wire  _T_3001;
  wire [6:0] _T_3007;
  wire [6:0] _T_3008;
  wire  _T_3010;
  wire [6:0] _T_3016;
  wire [6:0] _T_3017;
  wire  _T_3019;
  wire [6:0] _T_3025;
  wire [6:0] _T_3026;
  wire  _T_3028;
  wire [6:0] _T_3034;
  wire [6:0] _T_3035;
  wire  _T_3037;
  wire [6:0] _T_3043;
  wire [6:0] _T_3044;
  wire  _T_3046;
  wire [6:0] _T_3052;
  wire [6:0] _T_3053;
  wire  _T_3055;
  wire [6:0] _T_3061;
  wire [6:0] _T_3062;
  wire  _T_3064;
  wire [6:0] _T_3070;
  wire [6:0] _T_3071;
  wire  _T_3073;
  wire [6:0] _T_3079;
  wire [6:0] _T_3080;
  wire  _T_3082;
  wire [6:0] _T_3088;
  wire [6:0] _T_3089;
  wire  _T_3091;
  wire [6:0] _T_3097;
  wire [6:0] _T_3098;
  wire  _T_3100;
  wire [6:0] _T_3106;
  wire [6:0] _T_3107;
  wire  _T_3109;
  wire [6:0] _T_3115;
  wire [6:0] _T_3116;
  wire  _T_3118;
  wire [6:0] _T_3124;
  wire [6:0] _T_3125;
  wire  _T_3127;
  wire [6:0] _T_3133;
  wire [6:0] _T_3134;
  wire  _T_3136;
  wire [6:0] _T_3142;
  wire [6:0] _T_3143;
  wire  _T_3145;
  wire [6:0] _T_3151;
  wire [6:0] _T_3152;
  wire  _T_3154;
  wire [6:0] _T_3160;
  wire [6:0] _T_3161;
  wire  _T_3163;
  wire [6:0] _T_3169;
  wire [6:0] _T_3170;
  wire  _T_3172;
  wire  _T_3533;
  wire  _T_3534;
  wire  _T_3535;
  wire  _T_3536;
  wire [7:0] _T_3540;
  wire [7:0] _T_3544;
  wire [7:0] _T_3548;
  wire [7:0] _T_3552;
  wire [15:0] _T_3553;
  wire [15:0] _T_3554;
  wire [31:0] _T_3555;
  wire [7:0] _T_3579;
  wire  _T_3581;
  wire [7:0] _T_3583;
  wire  _T_3585;
  wire  _T_3594;
  wire  _T_3598;
  wire [7:0] _T_3599;
  wire [7:0] _GEN_60;
  wire [7:0] _T_3619;
  wire  _T_3621;
  wire [7:0] _T_3623;
  wire  _T_3625;
  wire  _T_3634;
  wire  _T_3638;
  wire [7:0] _T_3639;
  wire [7:0] _GEN_61;
  wire [15:0] _GEN_5671;
  wire [15:0] _T_3654;
  wire [15:0] _GEN_5672;
  wire [15:0] _T_3658;
  wire [7:0] _T_3659;
  wire  _T_3661;
  wire [7:0] _T_3663;
  wire  _T_3665;
  wire  _T_3674;
  wire  _T_3678;
  wire [7:0] _T_3679;
  wire [7:0] _GEN_62;
  wire [23:0] _GEN_5673;
  wire [23:0] _T_3694;
  wire [23:0] _GEN_5674;
  wire [23:0] _T_3698;
  wire [7:0] _T_3699;
  wire  _T_3701;
  wire [7:0] _T_3703;
  wire  _T_3705;
  wire  _T_3714;
  wire  _T_3718;
  wire [7:0] _T_3719;
  wire [7:0] _GEN_63;
  wire [31:0] _GEN_5675;
  wire [31:0] _T_3734;
  wire [31:0] _GEN_5676;
  wire [31:0] _T_3738;
  wire [31:0] _T_3743;
  wire  _T_3745;
  wire  _T_3758;
  wire [31:0] _GEN_64;
  wire  _T_3794;
  wire  _T_3798;
  wire [7:0] _GEN_65;
  wire  _T_3834;
  wire  _T_3838;
  wire [7:0] _GEN_66;
  wire [15:0] _GEN_5677;
  wire [15:0] _T_3854;
  wire [15:0] _GEN_5678;
  wire [15:0] _T_3858;
  wire  _T_3874;
  wire  _T_3878;
  wire [7:0] _GEN_67;
  wire [23:0] _GEN_5679;
  wire [23:0] _T_3894;
  wire [23:0] _GEN_5680;
  wire [23:0] _T_3898;
  wire  _T_3914;
  wire  _T_3918;
  wire [7:0] _GEN_68;
  wire [31:0] _GEN_5681;
  wire [31:0] _T_3934;
  wire [31:0] _GEN_5682;
  wire [31:0] _T_3938;
  wire  _T_3954;
  wire  _T_3958;
  wire [7:0] _GEN_69;
  wire  _T_3994;
  wire  _T_3998;
  wire [7:0] _GEN_70;
  wire [15:0] _GEN_5683;
  wire [15:0] _T_4014;
  wire [15:0] _GEN_5684;
  wire [15:0] _T_4018;
  wire  _T_4034;
  wire  _T_4038;
  wire [7:0] _GEN_71;
  wire [23:0] _GEN_5685;
  wire [23:0] _T_4054;
  wire [23:0] _GEN_5686;
  wire [23:0] _T_4058;
  wire  _T_4074;
  wire  _T_4078;
  wire [7:0] _GEN_72;
  wire [31:0] _GEN_5687;
  wire [31:0] _T_4094;
  wire [31:0] _GEN_5688;
  wire [31:0] _T_4098;
  wire  _T_4114;
  wire  _T_4118;
  wire [7:0] _GEN_73;
  wire  _T_4154;
  wire  _T_4158;
  wire [7:0] _GEN_74;
  wire [15:0] _GEN_5689;
  wire [15:0] _T_4174;
  wire [15:0] _GEN_5690;
  wire [15:0] _T_4178;
  wire  _T_4194;
  wire  _T_4198;
  wire [7:0] _GEN_75;
  wire [23:0] _GEN_5691;
  wire [23:0] _T_4214;
  wire [23:0] _GEN_5692;
  wire [23:0] _T_4218;
  wire  _T_4234;
  wire  _T_4238;
  wire [7:0] _GEN_76;
  wire [31:0] _GEN_5693;
  wire [31:0] _T_4254;
  wire [31:0] _GEN_5694;
  wire [31:0] _T_4258;
  wire  _T_4274;
  wire  _T_4278;
  wire [7:0] _GEN_77;
  wire  _T_4314;
  wire  _T_4318;
  wire [7:0] _GEN_78;
  wire [15:0] _GEN_5695;
  wire [15:0] _T_4334;
  wire [15:0] _GEN_5696;
  wire [15:0] _T_4338;
  wire  _T_4354;
  wire  _T_4358;
  wire [7:0] _GEN_79;
  wire [23:0] _GEN_5697;
  wire [23:0] _T_4374;
  wire [23:0] _GEN_5698;
  wire [23:0] _T_4378;
  wire  _T_4394;
  wire  _T_4398;
  wire [7:0] _GEN_80;
  wire [31:0] _GEN_5699;
  wire [31:0] _T_4414;
  wire [31:0] _GEN_5700;
  wire [31:0] _T_4418;
  wire  _T_4434;
  wire  _T_4438;
  wire [7:0] _GEN_81;
  wire  _T_4474;
  wire  _T_4478;
  wire [7:0] _GEN_82;
  wire [15:0] _GEN_5701;
  wire [15:0] _T_4494;
  wire [15:0] _GEN_5702;
  wire [15:0] _T_4498;
  wire  _T_4514;
  wire  _T_4518;
  wire [7:0] _GEN_83;
  wire [23:0] _GEN_5703;
  wire [23:0] _T_4534;
  wire [23:0] _GEN_5704;
  wire [23:0] _T_4538;
  wire  _T_4554;
  wire  _T_4558;
  wire [7:0] _GEN_84;
  wire [31:0] _GEN_5705;
  wire [31:0] _T_4574;
  wire [31:0] _GEN_5706;
  wire [31:0] _T_4578;
  wire  _T_4594;
  wire  _T_4598;
  wire [7:0] _GEN_85;
  wire  _T_4634;
  wire  _T_4638;
  wire [7:0] _GEN_86;
  wire [15:0] _GEN_5707;
  wire [15:0] _T_4654;
  wire [15:0] _GEN_5708;
  wire [15:0] _T_4658;
  wire  _T_4674;
  wire  _T_4678;
  wire [7:0] _GEN_87;
  wire [23:0] _GEN_5709;
  wire [23:0] _T_4694;
  wire [23:0] _GEN_5710;
  wire [23:0] _T_4698;
  wire  _T_4714;
  wire  _T_4718;
  wire [7:0] _GEN_88;
  wire [31:0] _GEN_5711;
  wire [31:0] _T_4734;
  wire [31:0] _GEN_5712;
  wire [31:0] _T_4738;
  wire  _T_4754;
  wire  _T_4758;
  wire [7:0] _GEN_89;
  wire  _T_4794;
  wire  _T_4798;
  wire [7:0] _GEN_90;
  wire [15:0] _GEN_5713;
  wire [15:0] _T_4814;
  wire [15:0] _GEN_5714;
  wire [15:0] _T_4818;
  wire  _T_4834;
  wire  _T_4838;
  wire [7:0] _GEN_91;
  wire [23:0] _GEN_5715;
  wire [23:0] _T_4854;
  wire [23:0] _GEN_5716;
  wire [23:0] _T_4858;
  wire  _T_4874;
  wire  _T_4878;
  wire [7:0] _GEN_92;
  wire [31:0] _GEN_5717;
  wire [31:0] _T_4894;
  wire [31:0] _GEN_5718;
  wire [31:0] _T_4898;
  wire  _T_4914;
  wire  _T_4918;
  wire [7:0] _GEN_93;
  wire  _T_4954;
  wire  _T_4958;
  wire [7:0] _GEN_94;
  wire [15:0] _GEN_5719;
  wire [15:0] _T_4974;
  wire [15:0] _GEN_5720;
  wire [15:0] _T_4978;
  wire  _T_4994;
  wire  _T_4998;
  wire [7:0] _GEN_95;
  wire [23:0] _GEN_5721;
  wire [23:0] _T_5014;
  wire [23:0] _GEN_5722;
  wire [23:0] _T_5018;
  wire  _T_5034;
  wire  _T_5038;
  wire [7:0] _GEN_96;
  wire [31:0] _GEN_5723;
  wire [31:0] _T_5054;
  wire [31:0] _GEN_5724;
  wire [31:0] _T_5058;
  wire  _T_5158;
  wire [31:0] _GEN_97;
  wire  _T_5194;
  wire  _T_5198;
  wire [7:0] _GEN_98;
  wire  _T_5234;
  wire  _T_5238;
  wire [7:0] _GEN_99;
  wire [15:0] _GEN_5725;
  wire [15:0] _T_5254;
  wire [15:0] _GEN_5726;
  wire [15:0] _T_5258;
  wire  _T_5274;
  wire  _T_5278;
  wire [7:0] _GEN_100;
  wire [23:0] _GEN_5727;
  wire [23:0] _T_5294;
  wire [23:0] _GEN_5728;
  wire [23:0] _T_5298;
  wire  _T_5314;
  wire  _T_5318;
  wire [7:0] _GEN_101;
  wire [31:0] _GEN_5729;
  wire [31:0] _T_5334;
  wire [31:0] _GEN_5730;
  wire [31:0] _T_5338;
  wire  _T_5354;
  wire  _T_5358;
  wire [7:0] _GEN_102;
  wire  _T_5394;
  wire  _T_5398;
  wire [7:0] _GEN_103;
  wire [15:0] _GEN_5731;
  wire [15:0] _T_5414;
  wire [15:0] _GEN_5732;
  wire [15:0] _T_5418;
  wire  _T_5434;
  wire  _T_5438;
  wire [7:0] _GEN_104;
  wire [23:0] _GEN_5733;
  wire [23:0] _T_5454;
  wire [23:0] _GEN_5734;
  wire [23:0] _T_5458;
  wire  _T_5474;
  wire  _T_5478;
  wire [7:0] _GEN_105;
  wire [31:0] _GEN_5735;
  wire [31:0] _T_5494;
  wire [31:0] _GEN_5736;
  wire [31:0] _T_5498;
  wire  _T_5514;
  wire  _T_5518;
  wire [7:0] _GEN_106;
  wire  _T_5554;
  wire  _T_5558;
  wire [7:0] _GEN_107;
  wire [15:0] _GEN_5737;
  wire [15:0] _T_5574;
  wire [15:0] _GEN_5738;
  wire [15:0] _T_5578;
  wire  _T_5594;
  wire  _T_5598;
  wire [7:0] _GEN_108;
  wire [23:0] _GEN_5739;
  wire [23:0] _T_5614;
  wire [23:0] _GEN_5740;
  wire [23:0] _T_5618;
  wire  _T_5634;
  wire  _T_5638;
  wire [7:0] _GEN_109;
  wire [31:0] _GEN_5741;
  wire [31:0] _T_5654;
  wire [31:0] _GEN_5742;
  wire [31:0] _T_5658;
  wire  _T_5714;
  wire  _T_5718;
  wire [7:0] _GEN_110;
  wire  _T_5754;
  wire  _T_5758;
  wire [7:0] _GEN_111;
  wire [15:0] _GEN_5743;
  wire [15:0] _T_5774;
  wire [15:0] _GEN_5744;
  wire [15:0] _T_5778;
  wire  _T_5794;
  wire  _T_5798;
  wire [7:0] _GEN_112;
  wire [23:0] _GEN_5745;
  wire [23:0] _T_5814;
  wire [23:0] _GEN_5746;
  wire [23:0] _T_5818;
  wire  _T_5834;
  wire  _T_5838;
  wire [7:0] _GEN_113;
  wire [31:0] _GEN_5747;
  wire [31:0] _T_5854;
  wire [31:0] _GEN_5748;
  wire [31:0] _T_5858;
  wire  _T_5874;
  wire  _T_5878;
  wire [7:0] _GEN_114;
  wire  _T_5914;
  wire  _T_5918;
  wire [7:0] _GEN_115;
  wire [15:0] _GEN_5749;
  wire [15:0] _T_5934;
  wire [15:0] _GEN_5750;
  wire [15:0] _T_5938;
  wire  _T_5954;
  wire  _T_5958;
  wire [7:0] _GEN_116;
  wire [23:0] _GEN_5751;
  wire [23:0] _T_5974;
  wire [23:0] _GEN_5752;
  wire [23:0] _T_5978;
  wire  _T_5994;
  wire  _T_5998;
  wire [7:0] _GEN_117;
  wire [31:0] _GEN_5753;
  wire [31:0] _T_6014;
  wire [31:0] _GEN_5754;
  wire [31:0] _T_6018;
  wire  _T_6038;
  wire [31:0] _GEN_118;
  wire  _T_6074;
  wire  _T_6078;
  wire [7:0] _GEN_119;
  wire  _T_6114;
  wire  _T_6118;
  wire [7:0] _GEN_120;
  wire [15:0] _GEN_5755;
  wire [15:0] _T_6134;
  wire [15:0] _GEN_5756;
  wire [15:0] _T_6138;
  wire  _T_6154;
  wire  _T_6158;
  wire [7:0] _GEN_121;
  wire [23:0] _GEN_5757;
  wire [23:0] _T_6174;
  wire [23:0] _GEN_5758;
  wire [23:0] _T_6178;
  wire  _T_6194;
  wire  _T_6198;
  wire [7:0] _GEN_122;
  wire [31:0] _GEN_5759;
  wire [31:0] _T_6214;
  wire [31:0] _GEN_5760;
  wire [31:0] _T_6218;
  wire  _T_6274;
  wire  _T_6278;
  wire [7:0] _GEN_123;
  wire  _T_6314;
  wire  _T_6318;
  wire [7:0] _GEN_124;
  wire [15:0] _GEN_5761;
  wire [15:0] _T_6334;
  wire [15:0] _GEN_5762;
  wire [15:0] _T_6338;
  wire  _T_6354;
  wire  _T_6358;
  wire [7:0] _GEN_125;
  wire [23:0] _GEN_5763;
  wire [23:0] _T_6374;
  wire [23:0] _GEN_5764;
  wire [23:0] _T_6378;
  wire  _T_6394;
  wire  _T_6398;
  wire [7:0] _GEN_126;
  wire [31:0] _GEN_5765;
  wire [31:0] _T_6414;
  wire [31:0] _GEN_5766;
  wire [31:0] _T_6418;
  wire  _T_6434;
  wire  _T_6438;
  wire [7:0] _GEN_127;
  wire  _T_6474;
  wire  _T_6478;
  wire [7:0] _GEN_128;
  wire [15:0] _GEN_5767;
  wire [15:0] _T_6494;
  wire [15:0] _GEN_5768;
  wire [15:0] _T_6498;
  wire  _T_6514;
  wire  _T_6518;
  wire [7:0] _GEN_129;
  wire [23:0] _GEN_5769;
  wire [23:0] _T_6534;
  wire [23:0] _GEN_5770;
  wire [23:0] _T_6538;
  wire  _T_6554;
  wire  _T_6558;
  wire [7:0] _GEN_130;
  wire [31:0] _GEN_5771;
  wire [31:0] _T_6574;
  wire [31:0] _GEN_5772;
  wire [31:0] _T_6578;
  wire  _T_6579;
  wire  _T_6580;
  wire  _T_6581;
  wire  _T_6582;
  wire  _T_6584;
  wire [1:0] _T_6586;
  wire [1:0] _T_6587;
  wire [2:0] _T_6588;
  wire [4:0] _T_6589;
  wire [31:0] _T_6602;
  wire  _T_6607;
  wire  _T_6609;
  wire  _T_6610;
  wire  _T_6611;
  wire  _T_6619;
  wire  _T_6620;
  wire  _T_6621;
  wire  _T_6622;
  wire  _T_6623;
  wire  _T_6624;
  wire  _T_6625;
  wire  _T_6626;
  wire  _T_6627;
  wire  _T_6628;
  wire  _T_6629;
  wire  _T_6630;
  wire  _T_6631;
  wire  _T_6632;
  wire  _T_6633;
  wire  _T_6634;
  wire  _T_6669;
  wire  _T_6670;
  wire  _T_6705;
  wire  _T_6801;
  wire  _T_6809;
  wire  _T_6817;
  wire  _T_6825;
  wire  _T_6833;
  wire  _T_6841;
  wire  _T_6849;
  wire  _T_6857;
  wire  _T_6865;
  wire  _T_6873;
  wire  _T_6881;
  wire  _T_6889;
  wire  _T_6897;
  wire  _T_6905;
  wire  _T_6913;
  wire  _T_6921;
  wire  _T_6966;
  wire  _T_6967;
  wire  _T_7002;
  wire  _T_7018;
  wire  _T_7026;
  wire  _T_7034;
  wire  _T_7098;
  wire  _T_7106;
  wire  _T_7114;
  wire  _T_7122;
  wire  _T_7130;
  wire  _T_7138;
  wire  _T_7146;
  wire  _T_7154;
  wire  _T_7162;
  wire  _T_7170;
  wire  _T_7178;
  wire  _T_7186;
  wire  _T_7194;
  wire  _T_7202;
  wire  _T_7210;
  wire  _T_7218;
  wire  _T_7298;
  wire  _T_7394;
  wire  _T_7402;
  wire  _T_7410;
  wire  _T_7418;
  wire  _T_7426;
  wire  _T_7434;
  wire  _T_7442;
  wire  _T_7450;
  wire  _T_7458;
  wire  _T_7466;
  wire  _T_7474;
  wire  _T_7482;
  wire  _T_7490;
  wire  _T_7498;
  wire  _T_7506;
  wire  _T_7514;
  wire  _T_7595;
  wire  _T_7611;
  wire  _T_7619;
  wire  _T_7627;
  wire  _T_7691;
  wire  _T_7699;
  wire  _T_7707;
  wire  _T_7715;
  wire  _T_7723;
  wire  _T_7731;
  wire  _T_7739;
  wire  _T_7747;
  wire  _T_7755;
  wire  _T_7763;
  wire  _T_7771;
  wire  _T_7779;
  wire  _T_7787;
  wire  _T_7795;
  wire  _T_7803;
  wire  _T_7811;
  wire  _GEN_255;
  wire  _GEN_256;
  wire  _GEN_257;
  wire  _GEN_258;
  wire  _GEN_259;
  wire  _GEN_260;
  wire  _GEN_261;
  wire  _GEN_262;
  wire  _GEN_263;
  wire  _GEN_264;
  wire  _GEN_265;
  wire  _GEN_266;
  wire  _GEN_267;
  wire  _GEN_268;
  wire  _GEN_269;
  wire  _GEN_270;
  wire  _GEN_271;
  wire  _GEN_272;
  wire  _GEN_273;
  wire  _GEN_274;
  wire  _GEN_275;
  wire  _GEN_276;
  wire  _GEN_277;
  wire  _GEN_278;
  wire  _GEN_279;
  wire  _GEN_280;
  wire  _GEN_281;
  wire  _GEN_282;
  wire  _GEN_283;
  wire  _GEN_284;
  wire  _GEN_285;
  wire [31:0] _GEN_286;
  wire [31:0] _GEN_287;
  wire [31:0] _GEN_288;
  wire [31:0] _GEN_289;
  wire [31:0] _GEN_290;
  wire [31:0] _GEN_291;
  wire [31:0] _GEN_292;
  wire [31:0] _GEN_293;
  wire [31:0] _GEN_294;
  wire [31:0] _GEN_295;
  wire [31:0] _GEN_296;
  wire [31:0] _GEN_297;
  wire [31:0] _GEN_298;
  wire [31:0] _GEN_299;
  wire [31:0] _GEN_300;
  wire [31:0] _GEN_301;
  wire [31:0] _GEN_302;
  wire [31:0] _GEN_303;
  wire [31:0] _GEN_304;
  wire [31:0] _GEN_305;
  wire [31:0] _GEN_306;
  wire [31:0] _GEN_307;
  wire [31:0] _GEN_308;
  wire [31:0] _GEN_309;
  wire [31:0] _GEN_310;
  wire [31:0] _GEN_311;
  wire [31:0] _GEN_312;
  wire [31:0] _GEN_313;
  wire [31:0] _GEN_314;
  wire [31:0] _GEN_315;
  wire [31:0] _GEN_316;
  wire [31:0] _T_7940;
  wire  _T_7941;
  wire [1:0] _T_7942;
  wire  _T_7956;
  wire [7:0] _GEN_317;
  wire  _T_7957;
  wire [7:0] _GEN_318;
  wire  _T_7958;
  wire [7:0] _GEN_319;
  wire  _T_7959;
  wire [7:0] _GEN_320;
  wire  _T_7960;
  wire [7:0] _GEN_321;
  wire  _T_7961;
  wire [7:0] _GEN_322;
  wire  _T_7962;
  wire [7:0] _GEN_323;
  wire  _T_7963;
  wire [7:0] _GEN_324;
  wire  _T_7964;
  wire [7:0] _GEN_325;
  wire  _T_7965;
  wire [7:0] _GEN_326;
  wire  _T_7966;
  wire [7:0] _GEN_327;
  wire  _T_7967;
  wire [7:0] _GEN_328;
  wire  _T_7968;
  wire [7:0] _GEN_329;
  wire  _T_7969;
  wire [7:0] _GEN_330;
  wire  _T_7970;
  wire [7:0] _GEN_331;
  wire  _T_7971;
  wire [7:0] _GEN_332;
  wire  _T_7972;
  wire [7:0] _GEN_333;
  wire  _T_7973;
  wire [7:0] _GEN_334;
  wire  _T_7974;
  wire [7:0] _GEN_335;
  wire  _T_7975;
  wire [7:0] _GEN_336;
  wire  _T_7976;
  wire [7:0] _GEN_337;
  wire  _T_7977;
  wire [7:0] _GEN_338;
  wire  _T_7978;
  wire [7:0] _GEN_339;
  wire  _T_7979;
  wire [7:0] _GEN_340;
  wire  _T_7980;
  wire [7:0] _GEN_341;
  wire  _T_7981;
  wire [7:0] _GEN_342;
  wire  _T_7982;
  wire [7:0] _GEN_343;
  wire  _T_7983;
  wire [7:0] _GEN_344;
  wire  _T_7984;
  wire [7:0] _GEN_345;
  wire  _T_7985;
  wire [7:0] _GEN_346;
  wire  _T_7986;
  wire [7:0] _GEN_347;
  wire  _T_7987;
  wire [7:0] _GEN_348;
  wire  _T_7988;
  wire [7:0] _GEN_349;
  wire  _T_7989;
  wire [7:0] _GEN_350;
  wire  _T_7990;
  wire [7:0] _GEN_351;
  wire  _T_7991;
  wire [7:0] _GEN_352;
  wire  _T_7992;
  wire [7:0] _GEN_353;
  wire  _T_7993;
  wire [7:0] _GEN_354;
  wire  _T_7994;
  wire [7:0] _GEN_355;
  wire  _T_7995;
  wire [7:0] _GEN_356;
  wire  _T_7996;
  wire [7:0] _GEN_357;
  wire  _T_7997;
  wire [7:0] _GEN_358;
  wire  _T_7998;
  wire [7:0] _GEN_359;
  wire  _T_7999;
  wire [7:0] _GEN_360;
  wire  _T_8000;
  wire [7:0] _GEN_361;
  wire  _T_8001;
  wire [7:0] _GEN_362;
  wire  _T_8002;
  wire [7:0] _GEN_363;
  wire  _T_8003;
  wire [7:0] _GEN_364;
  wire  _T_8004;
  wire [7:0] _GEN_365;
  wire  _T_8005;
  wire [7:0] _GEN_366;
  wire  _T_8006;
  wire [7:0] _GEN_367;
  wire  _T_8007;
  wire [7:0] _GEN_368;
  wire  _T_8008;
  wire [7:0] _GEN_369;
  wire  _T_8009;
  wire [7:0] _GEN_370;
  wire  _T_8010;
  wire [7:0] _GEN_371;
  wire  _T_8011;
  wire [7:0] _GEN_372;
  wire  _T_8012;
  wire [7:0] _GEN_373;
  wire  _T_8013;
  wire [7:0] _GEN_374;
  wire  _T_8014;
  wire [7:0] _GEN_375;
  wire  _T_8015;
  wire [7:0] _GEN_376;
  wire  _T_8016;
  wire [7:0] _GEN_377;
  wire  _T_8017;
  wire [7:0] _GEN_378;
  wire  _T_8018;
  wire [7:0] _GEN_379;
  wire  _T_8019;
  wire [7:0] _GEN_380;
  wire  _T_8020;
  wire [7:0] _GEN_381;
  wire  _T_8021;
  wire [7:0] _GEN_382;
  wire  _T_8022;
  wire [7:0] _GEN_383;
  wire  _T_8023;
  wire [7:0] _GEN_384;
  reg  goReg;
  reg [31:0] _RAND_83;
  wire  _GEN_385;
  wire  _GEN_386;
  wire  _T_8235;
  wire  _T_8236;
  wire  _T_8238;
  wire  _T_8239;
  wire  _T_8241;
  wire  _GEN_387;
  wire  _GEN_388;
  wire  _GEN_389;
  wire  _GEN_390;
  wire  _GEN_391;
  wire  _GEN_392;
  wire  _GEN_393;
  wire  _GEN_394;
  wire  _GEN_395;
  wire  _GEN_396;
  wire  _GEN_397;
  wire  _GEN_398;
  wire  _GEN_399;
  wire  _GEN_400;
  wire  _GEN_401;
  wire  _GEN_402;
  wire  _GEN_403;
  wire  _GEN_404;
  wire  _GEN_405;
  wire  _GEN_406;
  wire  _GEN_407;
  wire  _GEN_408;
  wire  _GEN_409;
  wire  _GEN_410;
  wire  _GEN_411;
  wire  _GEN_412;
  wire  _GEN_413;
  wire  _GEN_414;
  wire  _GEN_415;
  wire  _GEN_416;
  wire  _GEN_417;
  wire  _GEN_418;
  wire  _GEN_419;
  wire  _GEN_420;
  wire  _GEN_421;
  wire  _GEN_422;
  wire  _GEN_423;
  wire  _GEN_424;
  wire  _GEN_425;
  wire  _GEN_426;
  wire  _GEN_427;
  wire  _GEN_428;
  wire  _GEN_429;
  wire  _GEN_430;
  wire  _GEN_431;
  wire  _GEN_432;
  wire  _GEN_433;
  wire  _GEN_434;
  wire  _GEN_435;
  wire  _GEN_436;
  wire  _GEN_437;
  wire  _GEN_438;
  wire  _GEN_439;
  wire  _GEN_440;
  wire  _GEN_441;
  wire  _GEN_442;
  wire  _GEN_443;
  wire  _GEN_444;
  wire  _GEN_445;
  wire  _GEN_446;
  wire  _GEN_447;
  wire  _GEN_448;
  wire  _GEN_449;
  wire  _GEN_450;
  wire  _GEN_451;
  wire  _GEN_452;
  wire  _GEN_453;
  wire  _GEN_454;
  wire  _GEN_455;
  wire  _GEN_456;
  wire  _GEN_457;
  wire  _GEN_458;
  wire  _GEN_459;
  wire  _GEN_460;
  wire  _GEN_461;
  wire  _GEN_462;
  wire  _GEN_463;
  wire  _GEN_464;
  wire  _GEN_465;
  wire  _GEN_466;
  wire  _GEN_467;
  wire  _GEN_468;
  wire  _GEN_469;
  wire  _GEN_470;
  wire  _GEN_471;
  wire  _GEN_472;
  wire  _GEN_473;
  wire  _GEN_474;
  wire  _GEN_475;
  wire  _GEN_476;
  wire  _GEN_477;
  wire  _GEN_478;
  wire  _GEN_479;
  wire  _GEN_480;
  wire  _GEN_481;
  wire  _GEN_482;
  wire  _GEN_483;
  wire  _GEN_484;
  wire  _GEN_485;
  wire  _GEN_486;
  wire  _GEN_487;
  wire  _GEN_488;
  wire  _GEN_489;
  wire  _GEN_490;
  wire  _GEN_491;
  wire  _GEN_492;
  wire  _GEN_493;
  wire  _GEN_494;
  wire  _GEN_495;
  wire  _GEN_496;
  wire  _GEN_497;
  wire  _GEN_498;
  wire  _GEN_499;
  wire  _GEN_500;
  wire  _GEN_501;
  wire  _GEN_502;
  wire  _GEN_503;
  wire  _GEN_504;
  wire  _GEN_505;
  wire  _GEN_506;
  wire  _GEN_507;
  wire  _GEN_508;
  wire  _GEN_509;
  wire  _GEN_510;
  wire  _GEN_511;
  wire  _GEN_512;
  wire  _GEN_513;
  wire  _GEN_514;
  wire  _GEN_515;
  wire  _GEN_516;
  wire  _GEN_517;
  wire  _GEN_518;
  wire  _GEN_519;
  wire  _GEN_520;
  wire  _GEN_521;
  wire  _GEN_522;
  wire  _GEN_523;
  wire  _GEN_524;
  wire  _GEN_525;
  wire  _GEN_526;
  wire  _GEN_527;
  wire  _GEN_528;
  wire  _GEN_529;
  wire  _GEN_530;
  wire  _GEN_531;
  wire  _GEN_532;
  wire  _GEN_533;
  wire  _GEN_534;
  wire  _GEN_535;
  wire  _GEN_536;
  wire  _GEN_537;
  wire  _GEN_538;
  wire  _GEN_539;
  wire  _GEN_540;
  wire  _GEN_541;
  wire  _GEN_542;
  wire  _GEN_543;
  wire  _GEN_544;
  wire  _GEN_545;
  wire  _GEN_546;
  wire  _GEN_547;
  wire  _GEN_548;
  wire  _GEN_549;
  wire  _GEN_550;
  wire  _GEN_551;
  wire  _GEN_552;
  wire  _GEN_553;
  wire  _GEN_554;
  wire  _GEN_555;
  wire  _GEN_556;
  wire  _GEN_557;
  wire  _GEN_558;
  wire  _GEN_559;
  wire  _GEN_560;
  wire  _GEN_561;
  wire  _GEN_562;
  wire  _GEN_563;
  wire  _GEN_564;
  wire  _GEN_565;
  wire  _GEN_566;
  wire  _GEN_567;
  wire  _GEN_568;
  wire  _GEN_569;
  wire  _GEN_570;
  wire  _GEN_571;
  wire  _GEN_572;
  wire  _GEN_573;
  wire  _GEN_574;
  wire  _GEN_575;
  wire  _GEN_576;
  wire  _GEN_577;
  wire  _GEN_578;
  wire  _GEN_579;
  wire  _GEN_580;
  wire  _GEN_581;
  wire  _GEN_582;
  wire  _GEN_583;
  wire  _GEN_584;
  wire  _GEN_585;
  wire  _GEN_586;
  wire  _GEN_587;
  wire  _GEN_588;
  wire  _GEN_589;
  wire  _GEN_590;
  wire  _GEN_591;
  wire  _GEN_592;
  wire  _GEN_593;
  wire  _GEN_594;
  wire  _GEN_595;
  wire  _GEN_596;
  wire  _GEN_597;
  wire  _GEN_598;
  wire  _GEN_599;
  wire  _GEN_600;
  wire  _GEN_601;
  wire  _GEN_602;
  wire  _GEN_603;
  wire  _GEN_604;
  wire  _GEN_605;
  wire  _GEN_606;
  wire  _GEN_607;
  wire  _GEN_608;
  wire  _GEN_609;
  wire  _GEN_610;
  wire  _GEN_611;
  wire  _GEN_612;
  wire  _GEN_613;
  wire  _GEN_614;
  wire  _GEN_615;
  wire  _GEN_616;
  wire  _GEN_617;
  wire  _GEN_618;
  wire  _GEN_619;
  wire  _GEN_620;
  wire  _GEN_621;
  wire  _GEN_622;
  wire  _GEN_623;
  wire  _GEN_624;
  wire  _GEN_625;
  wire  _GEN_626;
  wire  _GEN_627;
  wire  _GEN_628;
  wire  _GEN_629;
  wire  _GEN_630;
  wire  _GEN_631;
  wire  _GEN_632;
  wire  _GEN_633;
  wire  _GEN_634;
  wire  _GEN_635;
  wire  _GEN_636;
  wire  _GEN_637;
  wire  _GEN_638;
  wire  _GEN_639;
  wire  _GEN_640;
  wire  _GEN_641;
  wire  _GEN_642;
  wire  _GEN_643;
  wire  _GEN_644;
  wire  _GEN_645;
  wire  _GEN_646;
  wire  _GEN_647;
  wire  _GEN_648;
  wire  _GEN_649;
  wire  _GEN_650;
  wire  _GEN_651;
  wire  _GEN_652;
  wire  _GEN_653;
  wire  _GEN_654;
  wire  _GEN_655;
  wire  _GEN_656;
  wire  _GEN_657;
  wire  _GEN_658;
  wire  _GEN_659;
  wire  _GEN_660;
  wire  _GEN_661;
  wire  _GEN_662;
  wire  _GEN_663;
  wire  _GEN_664;
  wire  _GEN_665;
  wire  _GEN_666;
  wire  _GEN_667;
  wire  _GEN_668;
  wire  _GEN_669;
  wire  _GEN_670;
  wire  _GEN_671;
  wire  _GEN_672;
  wire  _GEN_673;
  wire  _GEN_674;
  wire  _GEN_675;
  wire  _GEN_676;
  wire  _GEN_677;
  wire  _GEN_678;
  wire  _GEN_679;
  wire  _GEN_680;
  wire  _GEN_681;
  wire  _GEN_682;
  wire  _GEN_683;
  wire  _GEN_684;
  wire  _GEN_685;
  wire  _GEN_686;
  wire  _GEN_687;
  wire  _GEN_688;
  wire  _GEN_689;
  wire  _GEN_690;
  wire  _GEN_691;
  wire  _GEN_692;
  wire  _GEN_693;
  wire  _GEN_694;
  wire  _GEN_695;
  wire  _GEN_696;
  wire  _GEN_697;
  wire  _GEN_698;
  wire  _GEN_699;
  wire  _GEN_700;
  wire  _GEN_701;
  wire  _GEN_702;
  wire  _GEN_703;
  wire  _GEN_704;
  wire  _GEN_705;
  wire  _GEN_706;
  wire  _GEN_707;
  wire  _GEN_708;
  wire  _GEN_709;
  wire  _GEN_710;
  wire  _GEN_711;
  wire  _GEN_712;
  wire  _GEN_713;
  wire  _GEN_714;
  wire  _GEN_715;
  wire  _GEN_716;
  wire  _GEN_717;
  wire  _GEN_718;
  wire  _GEN_719;
  wire  _GEN_720;
  wire  _GEN_721;
  wire  _GEN_722;
  wire  _GEN_723;
  wire  _GEN_724;
  wire  _GEN_725;
  wire  _GEN_726;
  wire  _GEN_727;
  wire  _GEN_728;
  wire  _GEN_729;
  wire  _GEN_730;
  wire  _GEN_731;
  wire  _GEN_732;
  wire  _GEN_733;
  wire  _GEN_734;
  wire  _GEN_735;
  wire  _GEN_736;
  wire  _GEN_737;
  wire  _GEN_738;
  wire  _GEN_739;
  wire  _GEN_740;
  wire  _GEN_741;
  wire  _GEN_742;
  wire  _GEN_743;
  wire  _GEN_744;
  wire  _GEN_745;
  wire  _GEN_746;
  wire  _GEN_747;
  wire  _GEN_748;
  wire  _GEN_749;
  wire  _GEN_750;
  wire  _GEN_751;
  wire  _GEN_752;
  wire  _GEN_753;
  wire  _GEN_754;
  wire  _GEN_755;
  wire  _GEN_756;
  wire  _GEN_757;
  wire  _GEN_758;
  wire  _GEN_759;
  wire  _GEN_760;
  wire  _GEN_761;
  wire  _GEN_762;
  wire  _GEN_763;
  wire  _GEN_764;
  wire  _GEN_765;
  wire  _GEN_766;
  wire  _GEN_767;
  wire  _GEN_768;
  wire  _GEN_769;
  wire  _GEN_770;
  wire  _GEN_771;
  wire  _GEN_772;
  wire  _GEN_773;
  wire  _GEN_774;
  wire  _GEN_775;
  wire  _GEN_776;
  wire  _GEN_777;
  wire  _GEN_778;
  wire  _GEN_779;
  wire  _GEN_780;
  wire  _GEN_781;
  wire  _GEN_782;
  wire  _GEN_783;
  wire  _GEN_784;
  wire  _GEN_785;
  wire  _GEN_786;
  wire  _GEN_787;
  wire  _GEN_788;
  wire  _GEN_789;
  wire  _GEN_790;
  wire  _GEN_791;
  wire  _GEN_792;
  wire  _GEN_793;
  wire  _GEN_794;
  wire  _GEN_795;
  wire  _GEN_796;
  wire  _GEN_797;
  wire  _GEN_798;
  wire  _GEN_799;
  wire  _GEN_800;
  wire  _GEN_801;
  wire  _GEN_802;
  wire  _GEN_803;
  wire  _GEN_804;
  wire  _GEN_805;
  wire  _GEN_806;
  wire  _GEN_807;
  wire  _GEN_808;
  wire  _GEN_809;
  wire  _GEN_810;
  wire  _GEN_811;
  wire  _GEN_812;
  wire  _GEN_813;
  wire  _GEN_814;
  wire  _GEN_815;
  wire  _GEN_816;
  wire  _GEN_817;
  wire  _GEN_818;
  wire  _GEN_819;
  wire  _GEN_820;
  wire  _GEN_821;
  wire  _GEN_822;
  wire  _GEN_823;
  wire  _GEN_824;
  wire  _GEN_825;
  wire  _GEN_826;
  wire  _GEN_827;
  wire  _GEN_828;
  wire  _GEN_829;
  wire  _GEN_830;
  wire  _GEN_831;
  wire  _GEN_832;
  wire  _GEN_833;
  wire  _GEN_834;
  wire  _GEN_835;
  wire  _GEN_836;
  wire  _GEN_837;
  wire  _GEN_838;
  wire  _GEN_839;
  wire  _GEN_840;
  wire  _GEN_841;
  wire  _GEN_842;
  wire  _GEN_843;
  wire  _GEN_844;
  wire  _GEN_845;
  wire  _GEN_846;
  wire  _GEN_847;
  wire  _GEN_848;
  wire  _GEN_849;
  wire  _GEN_850;
  wire  _GEN_851;
  wire  _GEN_852;
  wire  _GEN_853;
  wire  _GEN_854;
  wire  _GEN_855;
  wire  _GEN_856;
  wire  _GEN_857;
  wire  _GEN_858;
  wire  _GEN_859;
  wire  _GEN_860;
  wire  _GEN_861;
  wire  _GEN_862;
  wire  _GEN_863;
  wire  _GEN_864;
  wire  _GEN_865;
  wire  _GEN_866;
  wire  _GEN_867;
  wire  _GEN_868;
  wire  _GEN_869;
  wire  _GEN_870;
  wire  _GEN_871;
  wire  _GEN_872;
  wire  _GEN_873;
  wire  _GEN_874;
  wire  _GEN_875;
  wire  _GEN_876;
  wire  _GEN_877;
  wire  _GEN_878;
  wire  _GEN_879;
  wire  _GEN_880;
  wire  _GEN_881;
  wire  _GEN_882;
  wire  _GEN_883;
  wire  _GEN_884;
  wire  _GEN_885;
  wire  _GEN_886;
  wire  _GEN_887;
  wire  _GEN_888;
  wire  _GEN_889;
  wire  _GEN_890;
  wire  _GEN_891;
  wire  _GEN_892;
  wire  _GEN_893;
  wire  _GEN_894;
  wire  _GEN_895;
  wire  _GEN_896;
  wire  _GEN_897;
  wire  _GEN_898;
  wire  _GEN_899;
  wire  _GEN_900;
  wire  _GEN_901;
  wire  _GEN_902;
  wire  _GEN_903;
  wire  _GEN_904;
  wire  _GEN_905;
  wire  _GEN_906;
  wire  _GEN_907;
  wire  _GEN_908;
  wire  _GEN_909;
  wire  _GEN_910;
  wire  _GEN_911;
  wire  _GEN_912;
  wire  _GEN_913;
  wire  _GEN_914;
  wire  _GEN_915;
  wire  _GEN_916;
  wire  _GEN_917;
  wire  _GEN_918;
  wire  _GEN_919;
  wire  _GEN_920;
  wire  _GEN_921;
  wire  _GEN_922;
  wire  _GEN_923;
  wire  _GEN_924;
  wire  _GEN_925;
  wire  _GEN_926;
  wire  _GEN_927;
  wire  _GEN_928;
  wire  _GEN_929;
  wire  _GEN_930;
  wire  _GEN_931;
  wire  _GEN_932;
  wire  _GEN_933;
  wire  _GEN_934;
  wire  _GEN_935;
  wire  _GEN_936;
  wire  _GEN_937;
  wire  _GEN_938;
  wire  _GEN_939;
  wire  _GEN_940;
  wire  _GEN_941;
  wire  _GEN_942;
  wire  _GEN_943;
  wire  _GEN_944;
  wire  _GEN_945;
  wire  _GEN_946;
  wire  _GEN_947;
  wire  _GEN_948;
  wire  _GEN_949;
  wire  _GEN_950;
  wire  _GEN_951;
  wire  _GEN_952;
  wire  _GEN_953;
  wire  _GEN_954;
  wire  _GEN_955;
  wire  _GEN_956;
  wire  _GEN_957;
  wire  _GEN_958;
  wire  _GEN_959;
  wire  _GEN_960;
  wire  _GEN_961;
  wire  _GEN_962;
  wire  _GEN_963;
  wire  _GEN_964;
  wire  _GEN_965;
  wire  _GEN_966;
  wire  _GEN_967;
  wire  _GEN_968;
  wire  _GEN_969;
  wire  _GEN_970;
  wire  _GEN_971;
  wire  _GEN_972;
  wire  _GEN_973;
  wire  _GEN_974;
  wire  _GEN_975;
  wire  _GEN_976;
  wire  _GEN_977;
  wire  _GEN_978;
  wire  _GEN_979;
  wire  _GEN_980;
  wire  _GEN_981;
  wire  _GEN_982;
  wire  _GEN_983;
  wire  _GEN_984;
  wire  _GEN_985;
  wire  _GEN_986;
  wire  _GEN_987;
  wire  _GEN_988;
  wire  _GEN_989;
  wire  _GEN_990;
  wire  _GEN_991;
  wire  _GEN_992;
  wire  _GEN_993;
  wire  _GEN_994;
  wire  _GEN_995;
  wire  _GEN_996;
  wire  _GEN_997;
  wire  _GEN_998;
  wire  _GEN_999;
  wire  _GEN_1000;
  wire  _GEN_1001;
  wire  _GEN_1002;
  wire  _GEN_1003;
  wire  _GEN_1004;
  wire  _GEN_1005;
  wire  _GEN_1006;
  wire  _GEN_1007;
  wire  _GEN_1008;
  wire  _GEN_1009;
  wire  _GEN_1010;
  wire  _GEN_1011;
  wire  _GEN_1012;
  wire  _GEN_1013;
  wire  _GEN_1014;
  wire  _GEN_1015;
  wire  _GEN_1016;
  wire  _GEN_1017;
  wire  _GEN_1018;
  wire  _GEN_1019;
  wire  _GEN_1020;
  wire  _GEN_1021;
  wire  _GEN_1022;
  wire  _GEN_1023;
  wire  _GEN_1024;
  wire  _GEN_1025;
  wire  _GEN_1026;
  wire  _GEN_1027;
  wire  _GEN_1028;
  wire  _GEN_1029;
  wire  _GEN_1030;
  wire  _GEN_1031;
  wire  _GEN_1032;
  wire  _GEN_1033;
  wire  _GEN_1034;
  wire  _GEN_1035;
  wire  _GEN_1036;
  wire  _GEN_1037;
  wire  _GEN_1038;
  wire  _GEN_1039;
  wire  _GEN_1040;
  wire  _GEN_1041;
  wire  _GEN_1042;
  wire  _GEN_1043;
  wire  _GEN_1044;
  wire  _GEN_1045;
  wire  _GEN_1046;
  wire  _GEN_1047;
  wire  _GEN_1048;
  wire  _GEN_1049;
  wire  _GEN_1050;
  wire  _GEN_1051;
  wire  _GEN_1052;
  wire  _GEN_1053;
  wire  _GEN_1054;
  wire  _GEN_1055;
  wire  _GEN_1056;
  wire  _GEN_1057;
  wire  _GEN_1058;
  wire  _GEN_1059;
  wire  _GEN_1060;
  wire  _GEN_1061;
  wire  _GEN_1062;
  wire  _GEN_1063;
  wire  _GEN_1064;
  wire  _GEN_1065;
  wire  _GEN_1066;
  wire  _GEN_1067;
  wire  _GEN_1068;
  wire  _GEN_1069;
  wire  _GEN_1070;
  wire  _GEN_1071;
  wire  _GEN_1072;
  wire  _GEN_1073;
  wire  _GEN_1074;
  wire  _GEN_1075;
  wire  _GEN_1076;
  wire  _GEN_1077;
  wire  _GEN_1078;
  wire  _GEN_1079;
  wire  _GEN_1080;
  wire  _GEN_1081;
  wire  _GEN_1082;
  wire  _GEN_1083;
  wire  _GEN_1084;
  wire  _GEN_1085;
  wire  _GEN_1086;
  wire  _GEN_1087;
  wire  _GEN_1088;
  wire  _GEN_1089;
  wire  _GEN_1090;
  wire  _GEN_1091;
  wire  _GEN_1092;
  wire  _GEN_1093;
  wire  _GEN_1094;
  wire  _GEN_1095;
  wire  _GEN_1096;
  wire  _GEN_1097;
  wire  _GEN_1098;
  wire  _GEN_1099;
  wire  _GEN_1100;
  wire  _GEN_1101;
  wire  _GEN_1102;
  wire  _GEN_1103;
  wire  _GEN_1104;
  wire  _GEN_1105;
  wire  _GEN_1106;
  wire  _GEN_1107;
  wire  _GEN_1108;
  wire  _GEN_1109;
  wire  _GEN_1110;
  wire  _GEN_1111;
  wire  _GEN_1112;
  wire  _GEN_1113;
  wire  _GEN_1114;
  wire  _GEN_1115;
  wire  _GEN_1116;
  wire  _GEN_1117;
  wire  _GEN_1118;
  wire  _GEN_1119;
  wire  _GEN_1120;
  wire  _GEN_1121;
  wire  _GEN_1122;
  wire  _GEN_1123;
  wire  _GEN_1124;
  wire  _GEN_1125;
  wire  _GEN_1126;
  wire  _GEN_1127;
  wire  _GEN_1128;
  wire  _GEN_1129;
  wire  _GEN_1130;
  wire  _GEN_1131;
  wire  _GEN_1132;
  wire  _GEN_1133;
  wire  _GEN_1134;
  wire  _GEN_1135;
  wire  _GEN_1136;
  wire  _GEN_1137;
  wire  _GEN_1138;
  wire  _GEN_1139;
  wire  _GEN_1140;
  wire  _GEN_1141;
  wire  _GEN_1142;
  wire  _GEN_1143;
  wire  _GEN_1144;
  wire  _GEN_1145;
  wire  _GEN_1146;
  wire  _GEN_1147;
  wire  _GEN_1148;
  wire  _GEN_1149;
  wire  _GEN_1150;
  wire  _GEN_1151;
  wire  _GEN_1152;
  wire  _GEN_1153;
  wire  _GEN_1154;
  wire  _GEN_1155;
  wire  _GEN_1156;
  wire  _GEN_1157;
  wire  _GEN_1158;
  wire  _GEN_1159;
  wire  _GEN_1160;
  wire  _GEN_1161;
  wire  _GEN_1162;
  wire  _GEN_1163;
  wire  _GEN_1164;
  wire  _GEN_1165;
  wire  _GEN_1166;
  wire  _GEN_1167;
  wire  _GEN_1168;
  wire  _GEN_1169;
  wire  _GEN_1170;
  wire  _GEN_1171;
  wire  _GEN_1172;
  wire  _GEN_1173;
  wire  _GEN_1174;
  wire  _GEN_1175;
  wire  _GEN_1176;
  wire  _GEN_1177;
  wire  _GEN_1178;
  wire  _GEN_1179;
  wire  _GEN_1180;
  wire  _GEN_1181;
  wire  _GEN_1182;
  wire  _GEN_1183;
  wire  _GEN_1184;
  wire  _GEN_1185;
  wire  _GEN_1186;
  wire  _GEN_1187;
  wire  _GEN_1188;
  wire  _GEN_1189;
  wire  _GEN_1190;
  wire  _GEN_1191;
  wire  _GEN_1192;
  wire  _GEN_1193;
  wire  _GEN_1194;
  wire  _GEN_1195;
  wire  _GEN_1196;
  wire  _GEN_1197;
  wire  _GEN_1198;
  wire  _GEN_1199;
  wire  _GEN_1200;
  wire  _GEN_1201;
  wire  _GEN_1202;
  wire  _GEN_1203;
  wire  _GEN_1204;
  wire  _GEN_1205;
  wire  _GEN_1206;
  wire  _GEN_1207;
  wire  _GEN_1208;
  wire  _GEN_1209;
  wire  _GEN_1210;
  wire  _GEN_1211;
  wire  _GEN_1212;
  wire  _GEN_1213;
  wire  _GEN_1214;
  wire  _GEN_1215;
  wire  _GEN_1216;
  wire  _GEN_1217;
  wire  _GEN_1218;
  wire  _GEN_1219;
  wire  _GEN_1220;
  wire  _GEN_1221;
  wire  _GEN_1222;
  wire  _GEN_1223;
  wire  _GEN_1224;
  wire  _GEN_1225;
  wire  _GEN_1226;
  wire  _GEN_1227;
  wire  _GEN_1228;
  wire  _GEN_1229;
  wire  _GEN_1230;
  wire  _GEN_1231;
  wire  _GEN_1232;
  wire  _GEN_1233;
  wire  _GEN_1234;
  wire  _GEN_1235;
  wire  _GEN_1236;
  wire  _GEN_1237;
  wire  _GEN_1238;
  wire  _GEN_1239;
  wire  _GEN_1240;
  wire  _GEN_1241;
  wire  _GEN_1242;
  wire  _GEN_1243;
  wire  _GEN_1244;
  wire  _GEN_1245;
  wire  _GEN_1246;
  wire  _GEN_1247;
  wire  _GEN_1248;
  wire  _GEN_1249;
  wire  _GEN_1250;
  wire  _GEN_1251;
  wire  _GEN_1252;
  wire  _GEN_1253;
  wire  _GEN_1254;
  wire  _GEN_1255;
  wire  _GEN_1256;
  wire  _GEN_1257;
  wire  _GEN_1258;
  wire  _GEN_1259;
  wire  _GEN_1260;
  wire  _GEN_1261;
  wire  _GEN_1262;
  wire  _GEN_1263;
  wire  _GEN_1264;
  wire  _GEN_1265;
  wire  _GEN_1266;
  wire  _GEN_1267;
  wire  _GEN_1268;
  wire  _GEN_1269;
  wire  _GEN_1270;
  wire  _GEN_1271;
  wire  _GEN_1272;
  wire  _GEN_1273;
  wire  _GEN_1274;
  wire  _GEN_1275;
  wire  _GEN_1276;
  wire  _GEN_1277;
  wire  _GEN_1278;
  wire  _GEN_1279;
  wire  _GEN_1280;
  wire  _GEN_1281;
  wire  _GEN_1282;
  wire  _GEN_1283;
  wire  _GEN_1284;
  wire  _GEN_1285;
  wire  _GEN_1286;
  wire  _GEN_1287;
  wire  _GEN_1288;
  wire  _GEN_1289;
  wire  _GEN_1290;
  wire  _GEN_1291;
  wire  _GEN_1292;
  wire  _GEN_1293;
  wire  _GEN_1294;
  wire  _GEN_1295;
  wire  _GEN_1296;
  wire  _GEN_1297;
  wire  _GEN_1298;
  wire  _GEN_1299;
  wire  _GEN_1300;
  wire  _GEN_1301;
  wire  _GEN_1302;
  wire  _GEN_1303;
  wire  _GEN_1304;
  wire  _GEN_1305;
  wire  _GEN_1306;
  wire  _GEN_1307;
  wire  _GEN_1308;
  wire  _GEN_1309;
  wire  _GEN_1310;
  wire  _GEN_1311;
  wire  _GEN_1312;
  wire  _GEN_1313;
  wire  _GEN_1314;
  wire  _GEN_1315;
  wire  _GEN_1316;
  wire  _GEN_1317;
  wire  _GEN_1318;
  wire  _GEN_1319;
  wire  _GEN_1320;
  wire  _GEN_1321;
  wire  _GEN_1322;
  wire  _GEN_1323;
  wire  _GEN_1324;
  wire  _GEN_1325;
  wire  _GEN_1326;
  wire  _GEN_1327;
  wire  _GEN_1328;
  wire  _GEN_1329;
  wire  _GEN_1330;
  wire  _GEN_1331;
  wire  _GEN_1332;
  wire  _GEN_1333;
  wire  _GEN_1334;
  wire  _GEN_1335;
  wire  _GEN_1336;
  wire  _GEN_1337;
  wire  _GEN_1338;
  wire  _GEN_1339;
  wire  _GEN_1340;
  wire  _GEN_1341;
  wire  _GEN_1342;
  wire  _GEN_1343;
  wire  _GEN_1344;
  wire  _GEN_1345;
  wire  _GEN_1346;
  wire  _GEN_1347;
  wire  _GEN_1348;
  wire  _GEN_1349;
  wire  _GEN_1350;
  wire  _GEN_1351;
  wire  _GEN_1352;
  wire  _GEN_1353;
  wire  _GEN_1354;
  wire  _GEN_1355;
  wire  _GEN_1356;
  wire  _GEN_1357;
  wire  _GEN_1358;
  wire  _GEN_1359;
  wire  _GEN_1360;
  wire  _GEN_1361;
  wire  _GEN_1362;
  wire  _GEN_1363;
  wire  _GEN_1364;
  wire  _GEN_1365;
  wire  _GEN_1366;
  wire  _GEN_1367;
  wire  _GEN_1368;
  wire  _GEN_1369;
  wire  _GEN_1370;
  wire  _GEN_1371;
  wire  _GEN_1372;
  wire  _GEN_1373;
  wire  _GEN_1374;
  wire  _GEN_1375;
  wire  _GEN_1376;
  wire  _GEN_1377;
  wire  _GEN_1378;
  wire  _GEN_1379;
  wire  _GEN_1380;
  wire  _GEN_1381;
  wire  _GEN_1382;
  wire  _GEN_1383;
  wire  _GEN_1384;
  wire  _GEN_1385;
  wire  _GEN_1386;
  wire  _GEN_1387;
  wire  _GEN_1388;
  wire  _GEN_1389;
  wire  _GEN_1390;
  wire  _GEN_1391;
  wire  _GEN_1392;
  wire  _GEN_1393;
  wire  _GEN_1394;
  wire  _GEN_1395;
  wire  _GEN_1396;
  wire  _GEN_1397;
  wire  _GEN_1398;
  wire  _GEN_1399;
  wire  _GEN_1400;
  wire  _GEN_1401;
  wire  _GEN_1402;
  wire  _GEN_1403;
  wire  _GEN_1404;
  wire  _GEN_1405;
  wire  _GEN_1406;
  wire  _GEN_1407;
  wire  _GEN_1408;
  wire  _GEN_1409;
  wire  _GEN_1410;
  wire  _GEN_1411;
  wire  _GEN_1412;
  wire [15:0] _T_23654;
  wire  _T_23655;
  wire  _T_23656;
  wire  _T_23657;
  wire [2:0] _T_23659;
  reg [31:0] abstractGeneratedMem_0;
  reg [31:0] _RAND_84;
  reg [31:0] abstractGeneratedMem_1;
  reg [31:0] _RAND_85;
  wire [4:0] abstractGeneratedI_rd;
  wire [4:0] abstractGeneratedS_rs2;
  wire [15:0] _T_23685;
  wire [11:0] _T_23719;
  wire [19:0] _T_23721;
  wire [31:0] _T_23722;
  wire [7:0] _T_23723;
  wire [14:0] _T_23724;
  wire [11:0] _T_23725;
  wire [16:0] _T_23726;
  wire [31:0] _T_23727;
  wire [31:0] _T_23728;
  wire [31:0] _T_23733;
  wire [31:0] _T_23739;
  wire [31:0] _GEN_2437;
  wire [31:0] _GEN_2438;
  wire [6:0] _T_23745;
  wire [7:0] _T_23746;
  wire [7:0] _T_23748;
  wire [7:0] _T_23750;
  wire [7:0] _T_23752;
  wire [7:0] _T_23754;
  wire [7:0] _T_23756;
  wire [7:0] _T_23758;
  wire [7:0] _T_23760;
  wire [7:0] _T_23762;
  wire [7:0] _T_23764;
  wire [7:0] _T_23766;
  wire [7:0] _T_23768;
  wire [7:0] _T_23770;
  wire [7:0] _T_23772;
  wire [7:0] _T_23774;
  wire [7:0] _T_23776;
  wire [7:0] _T_23778;
  wire [7:0] _T_23780;
  wire [7:0] _T_23782;
  wire [7:0] _T_23784;
  wire [7:0] _T_23786;
  wire [7:0] _T_23788;
  wire [7:0] _T_23790;
  wire [7:0] _T_23792;
  wire [7:0] _T_23794;
  wire [7:0] _T_23796;
  wire [7:0] _T_23798;
  wire [7:0] _T_23800;
  wire [7:0] _T_23802;
  wire [7:0] _T_23804;
  wire [7:0] _T_23806;
  wire [7:0] _T_23808;
  wire [7:0] _T_23810;
  wire [7:0] _T_23812;
  wire [7:0] _T_23814;
  wire [7:0] _T_23816;
  wire [7:0] _T_23818;
  wire [7:0] _T_23820;
  wire [7:0] _T_23822;
  wire [7:0] _T_23824;
  wire [7:0] _T_23826;
  wire [7:0] _T_23828;
  wire [7:0] _T_23830;
  wire [7:0] _T_23832;
  wire [7:0] _T_23834;
  wire [7:0] _T_23836;
  wire [7:0] _T_23838;
  wire [7:0] _T_23840;
  wire [7:0] _T_23842;
  wire [7:0] _T_23844;
  wire [7:0] _T_23846;
  wire [7:0] _T_23848;
  wire [7:0] _T_23850;
  wire [7:0] _T_23852;
  wire [7:0] _T_23854;
  wire [7:0] _T_23856;
  wire [7:0] _T_23858;
  wire [7:0] _T_23860;
  wire [7:0] _T_23862;
  wire [7:0] _T_23864;
  wire [7:0] _T_23866;
  wire [7:0] _T_23868;
  wire [7:0] _T_23870;
  wire [7:0] _T_23872;
  wire [7:0] _T_23874;
  wire [7:0] _T_23876;
  wire [7:0] _T_23878;
  wire [7:0] _T_23880;
  wire [7:0] _T_23882;
  wire [7:0] _T_23884;
  wire [7:0] _T_23886;
  wire [7:0] _T_23888;
  wire [7:0] _T_23890;
  wire [7:0] _T_23892;
  wire [7:0] _T_23894;
  wire [7:0] _T_23896;
  wire [7:0] _T_23898;
  wire [7:0] _T_23900;
  wire [7:0] _T_23902;
  wire [7:0] _T_23904;
  wire [7:0] _T_23906;
  wire [7:0] _T_23908;
  wire [7:0] _T_23910;
  wire [7:0] _T_23912;
  wire [7:0] _T_23914;
  wire [7:0] _T_23916;
  wire [7:0] _T_23918;
  wire [7:0] _T_23920;
  wire [7:0] _T_23922;
  wire [7:0] _T_23924;
  wire [7:0] _T_23926;
  wire [7:0] _T_23928;
  wire [7:0] _T_23930;
  wire [7:0] _T_23932;
  wire [7:0] _T_23934;
  wire [7:0] _T_23936;
  wire [7:0] _T_23938;
  wire [7:0] _T_23940;
  wire [7:0] _T_23942;
  wire [7:0] _T_23944;
  wire [7:0] _T_23946;
  wire [7:0] _T_23948;
  wire [7:0] _T_23950;
  wire [7:0] _T_23952;
  wire [7:0] _T_23954;
  wire [7:0] _T_23956;
  wire [7:0] _T_23958;
  wire [7:0] _T_23960;
  wire [7:0] _T_23962;
  wire [7:0] _T_23964;
  wire [7:0] _T_23966;
  wire [7:0] _T_23968;
  wire [7:0] _T_23970;
  wire [7:0] _T_23972;
  wire [7:0] _T_23974;
  wire [7:0] _T_23976;
  wire [7:0] _T_23978;
  wire [7:0] _T_23980;
  wire [7:0] _T_23982;
  wire [7:0] _T_23984;
  wire [7:0] _T_23986;
  wire [7:0] _T_23988;
  wire [7:0] _T_23990;
  wire [7:0] _T_23992;
  wire [7:0] _T_23994;
  wire [7:0] _T_23996;
  wire [7:0] _T_23998;
  wire [7:0] _T_24000;
  wire [7:0] _T_24002;
  wire [7:0] _T_24004;
  wire [7:0] _T_24006;
  wire [7:0] _T_24008;
  wire [7:0] _T_24010;
  wire [7:0] _T_24012;
  wire [7:0] _T_24014;
  wire [7:0] _T_24016;
  wire [7:0] _T_24018;
  wire [7:0] _T_24020;
  wire [7:0] _T_24022;
  wire [7:0] _T_24024;
  wire [7:0] _T_24026;
  wire [7:0] _T_24028;
  wire [7:0] _T_24030;
  wire [7:0] _T_24032;
  wire [7:0] _T_24034;
  wire [7:0] _T_24036;
  wire [7:0] _T_24038;
  wire [7:0] _T_24040;
  wire [7:0] _T_24042;
  wire [7:0] _T_24044;
  wire [7:0] _T_24046;
  wire [7:0] _T_24048;
  wire [7:0] _T_24050;
  wire [7:0] _T_24052;
  wire [7:0] _T_24054;
  wire [7:0] _T_24056;
  wire [7:0] _T_24058;
  wire [7:0] _T_24060;
  wire [7:0] _T_24062;
  wire [7:0] _T_24064;
  wire [7:0] _T_24066;
  wire [7:0] _T_24068;
  wire [7:0] _T_24070;
  wire [7:0] _T_24072;
  wire [7:0] _T_24074;
  wire [7:0] _T_24076;
  wire [7:0] _T_24078;
  wire [7:0] _T_24080;
  wire [7:0] _T_24082;
  wire [7:0] _T_24084;
  wire [7:0] _T_24086;
  wire [7:0] _T_24088;
  wire [7:0] _T_24090;
  wire [7:0] _T_24092;
  wire [7:0] _T_24094;
  wire [7:0] _T_24096;
  wire [7:0] _T_24098;
  wire [7:0] _T_24100;
  wire [7:0] _T_24102;
  wire [7:0] _T_24104;
  wire [7:0] _T_24106;
  wire [7:0] _T_24108;
  wire [7:0] _T_24110;
  wire [7:0] _T_24112;
  wire [7:0] _T_24114;
  wire [7:0] _T_24116;
  wire [7:0] _T_24118;
  wire [7:0] _T_24120;
  wire [7:0] _T_24122;
  wire [7:0] _T_24124;
  wire [7:0] _T_24126;
  wire [7:0] _T_24128;
  wire [7:0] _T_24130;
  wire [7:0] _T_24132;
  wire [7:0] _T_24134;
  wire [7:0] _T_24136;
  wire [7:0] _T_24138;
  wire [7:0] _T_24140;
  wire [7:0] _T_24142;
  wire [7:0] _T_24144;
  wire [7:0] _T_24146;
  wire [7:0] _T_24148;
  wire [7:0] _T_24150;
  wire [7:0] _T_24152;
  wire [7:0] _T_24154;
  wire [7:0] _T_24156;
  wire [7:0] _T_24158;
  wire [7:0] _T_24160;
  wire [7:0] _T_24162;
  wire [7:0] _T_24164;
  wire [7:0] _T_24166;
  wire [7:0] _T_24168;
  wire [7:0] _T_24170;
  wire [7:0] _T_24172;
  wire [7:0] _T_24174;
  wire [7:0] _T_24176;
  wire [7:0] _T_24178;
  wire [7:0] _T_24180;
  wire [7:0] _T_24182;
  wire [7:0] _T_24184;
  wire [7:0] _T_24186;
  wire [7:0] _T_24188;
  wire [7:0] _T_24190;
  wire [7:0] _T_24192;
  wire [7:0] _T_24194;
  wire [7:0] _T_24196;
  wire [7:0] _T_24198;
  wire [7:0] _T_24200;
  wire [7:0] _T_24202;
  wire [7:0] _T_24204;
  wire [7:0] _T_24206;
  wire [7:0] _T_24208;
  wire [7:0] _T_24210;
  wire [7:0] _T_24212;
  wire [7:0] _T_24214;
  wire [7:0] _T_24216;
  wire [7:0] _T_24218;
  wire [7:0] _T_24220;
  wire [7:0] _T_24222;
  wire [7:0] _T_24224;
  wire [7:0] _T_24226;
  wire [7:0] _T_24228;
  wire [7:0] _T_24230;
  wire [7:0] _T_24232;
  wire [7:0] _T_24234;
  wire [7:0] _T_24236;
  wire [7:0] _T_24238;
  wire [7:0] _T_24240;
  wire [7:0] _T_24242;
  wire [7:0] _T_24244;
  wire [7:0] _T_24246;
  wire [7:0] _T_24248;
  wire [7:0] _T_24250;
  wire [7:0] _T_24252;
  wire [7:0] _T_24254;
  wire [7:0] _T_24256;
  wire [7:0] _T_24258;
  wire [7:0] _T_24260;
  wire [7:0] _T_24262;
  wire [7:0] _T_24264;
  wire [7:0] _T_24266;
  wire [7:0] _T_24268;
  wire [7:0] _T_24270;
  wire [7:0] _T_24272;
  wire [7:0] _T_24274;
  wire [7:0] _T_24276;
  wire [7:0] _T_24278;
  wire [7:0] _T_24280;
  wire [7:0] _T_24282;
  wire [7:0] _T_24284;
  wire [7:0] _T_24286;
  wire [7:0] _T_24288;
  wire [7:0] _T_24290;
  wire [7:0] _T_24292;
  wire [7:0] _T_24294;
  wire [7:0] _T_24296;
  wire [7:0] _T_24298;
  wire [7:0] _T_24300;
  wire [7:0] _T_24302;
  wire [7:0] _T_24304;
  wire [7:0] _T_24306;
  wire [7:0] _T_24308;
  wire [7:0] _T_24310;
  wire [7:0] _T_24312;
  wire [7:0] _T_24314;
  wire [7:0] _T_24316;
  wire [7:0] _T_24318;
  wire [7:0] _T_24320;
  wire [7:0] _T_24322;
  wire [7:0] _T_24324;
  wire [7:0] _T_24326;
  wire [7:0] _T_24328;
  wire [7:0] _T_24330;
  wire [7:0] _T_24332;
  wire [7:0] _T_24334;
  wire [7:0] _T_24336;
  wire [7:0] _T_24338;
  wire [7:0] _T_24340;
  wire [7:0] _T_24342;
  wire [7:0] _T_24344;
  wire [7:0] _T_24346;
  wire [7:0] _T_24348;
  wire [7:0] _T_24350;
  wire [7:0] _T_24352;
  wire [7:0] _T_24354;
  wire [7:0] _T_24356;
  wire [7:0] _T_24358;
  wire [7:0] _T_24360;
  wire [7:0] _T_24362;
  wire [7:0] _T_24364;
  wire [7:0] _T_24366;
  wire [7:0] _T_24368;
  wire [7:0] _T_24370;
  wire [7:0] _T_24372;
  wire [7:0] _T_24374;
  wire [7:0] _T_24376;
  wire [7:0] _T_24378;
  wire [7:0] _T_24380;
  wire [7:0] _T_24382;
  wire [7:0] _T_24384;
  wire [7:0] _T_24386;
  wire [7:0] _T_24388;
  wire [7:0] _T_24390;
  wire [7:0] _T_24392;
  wire [7:0] _T_24394;
  wire [7:0] _T_24396;
  wire [7:0] _T_24398;
  wire [7:0] _T_24400;
  wire [7:0] _T_24402;
  wire [7:0] _T_24404;
  wire [7:0] _T_24406;
  wire [7:0] _T_24408;
  wire [7:0] _T_24410;
  wire [7:0] _T_24412;
  wire [7:0] _T_24414;
  wire [7:0] _T_24416;
  wire [7:0] _T_24418;
  wire [7:0] _T_24420;
  wire [7:0] _T_24422;
  wire [7:0] _T_24424;
  wire [7:0] _T_24426;
  wire [7:0] _T_24428;
  wire [7:0] _T_24430;
  wire [7:0] _T_24432;
  wire [7:0] _T_24434;
  wire [7:0] _T_24436;
  wire [7:0] _T_24438;
  wire [7:0] _T_24440;
  wire [7:0] _T_24442;
  wire [7:0] _T_24444;
  wire [7:0] _T_24446;
  wire [7:0] _T_24448;
  wire [7:0] _T_24450;
  wire [7:0] _T_24452;
  wire [7:0] _T_24454;
  wire [7:0] _T_24456;
  wire [7:0] _T_24458;
  wire [7:0] _T_24460;
  wire [7:0] _T_24462;
  wire [7:0] _T_24464;
  wire [7:0] _T_24466;
  wire [7:0] _T_24468;
  wire [7:0] _T_24470;
  wire [7:0] _T_24472;
  wire [7:0] _T_24474;
  wire [7:0] _T_24476;
  wire [7:0] _T_24478;
  wire [7:0] _T_24480;
  wire [7:0] _T_24482;
  wire [7:0] _T_24484;
  wire [7:0] _T_24486;
  wire [7:0] _T_24488;
  wire [7:0] _T_24490;
  wire [7:0] _T_24492;
  wire [7:0] _T_24494;
  wire [7:0] _T_24496;
  wire [7:0] _T_24498;
  wire [7:0] _T_24500;
  wire [7:0] _T_24502;
  wire [7:0] _T_24504;
  wire [7:0] _T_24506;
  wire [7:0] _T_24508;
  wire [7:0] _T_24510;
  wire [7:0] _T_24512;
  wire [7:0] _T_24514;
  wire [7:0] _T_24516;
  wire [7:0] _T_24518;
  wire [7:0] _T_24520;
  wire [7:0] _T_24522;
  wire [7:0] _T_24524;
  wire [7:0] _T_24526;
  wire [7:0] _T_24528;
  wire [7:0] _T_24530;
  wire [7:0] _T_24532;
  wire [7:0] _T_24534;
  wire [7:0] _T_24536;
  wire [7:0] _T_24538;
  wire [7:0] _T_24540;
  wire [7:0] _T_24542;
  wire [7:0] _T_24544;
  wire [7:0] _T_24546;
  wire [7:0] _T_24548;
  wire [7:0] _T_24550;
  wire [7:0] _T_24552;
  wire [7:0] _T_24554;
  wire [7:0] _T_24556;
  wire [7:0] _T_24558;
  wire [7:0] _T_24560;
  wire [7:0] _T_24562;
  wire [7:0] _T_24564;
  wire [7:0] _T_24566;
  wire [7:0] _T_24568;
  wire [7:0] _T_24570;
  wire [7:0] _T_24572;
  wire [7:0] _T_24574;
  wire [7:0] _T_24576;
  wire [7:0] _T_24578;
  wire [7:0] _T_24580;
  wire [7:0] _T_24582;
  wire [7:0] _T_24584;
  wire [7:0] _T_24586;
  wire [7:0] _T_24588;
  wire [7:0] _T_24590;
  wire [7:0] _T_24592;
  wire [7:0] _T_24594;
  wire [7:0] _T_24596;
  wire [7:0] _T_24598;
  wire [7:0] _T_24600;
  wire [7:0] _T_24602;
  wire [7:0] _T_24604;
  wire [7:0] _T_24606;
  wire [7:0] _T_24608;
  wire [7:0] _T_24610;
  wire [7:0] _T_24612;
  wire [7:0] _T_24614;
  wire [7:0] _T_24616;
  wire [7:0] _T_24618;
  wire [7:0] _T_24620;
  wire [7:0] _T_24622;
  wire [7:0] _T_24624;
  wire [7:0] _T_24626;
  wire [7:0] _T_24628;
  wire [7:0] _T_24630;
  wire [7:0] _T_24632;
  wire [7:0] _T_24634;
  wire [7:0] _T_24636;
  wire [7:0] _T_24638;
  wire [7:0] _T_24640;
  wire [7:0] _T_24642;
  wire [7:0] _T_24644;
  wire [7:0] _T_24646;
  wire [7:0] _T_24648;
  wire [7:0] _T_24650;
  wire [7:0] _T_24652;
  wire [7:0] _T_24654;
  wire [7:0] _T_24656;
  wire [7:0] _T_24658;
  wire [7:0] _T_24660;
  wire [7:0] _T_24662;
  wire [7:0] _T_24664;
  wire [7:0] _T_24666;
  wire [7:0] _T_24668;
  wire [7:0] _T_24670;
  wire [7:0] _T_24672;
  wire [7:0] _T_24674;
  wire [7:0] _T_24676;
  wire [7:0] _T_24678;
  wire [7:0] _T_24680;
  wire [7:0] _T_24682;
  wire [7:0] _T_24684;
  wire [7:0] _T_24686;
  wire [7:0] _T_24688;
  wire [7:0] _T_24690;
  wire [7:0] _T_24692;
  wire [7:0] _T_24694;
  wire [7:0] _T_24696;
  wire [7:0] _T_24698;
  wire [7:0] _T_24700;
  wire [7:0] _T_24702;
  wire [7:0] _T_24704;
  wire [7:0] _T_24706;
  wire [7:0] _T_24708;
  wire [7:0] _T_24710;
  wire [7:0] _T_24712;
  wire [7:0] _T_24714;
  wire [7:0] _T_24716;
  wire [7:0] _T_24718;
  wire [7:0] _T_24720;
  wire [7:0] _T_24722;
  wire [7:0] _T_24724;
  wire [7:0] _T_24726;
  wire [7:0] _T_24728;
  wire [7:0] _T_24730;
  wire [7:0] _T_24732;
  wire [7:0] _T_24734;
  wire [7:0] _T_24736;
  wire [7:0] _T_24738;
  wire [7:0] _T_24740;
  wire [7:0] _T_24742;
  wire [7:0] _T_24744;
  wire [7:0] _T_24746;
  wire [7:0] _T_24748;
  wire [7:0] _T_24750;
  wire [7:0] _T_24752;
  wire [7:0] _T_24754;
  wire [7:0] _T_24756;
  wire [7:0] _T_24758;
  wire [7:0] _T_24760;
  wire [7:0] _T_24762;
  wire [7:0] _T_24764;
  wire [7:0] _T_24766;
  wire [7:0] _T_24768;
  wire [7:0] _T_24770;
  wire [7:0] _T_24772;
  wire [7:0] _T_24774;
  wire [7:0] _T_24776;
  wire [7:0] _T_24778;
  wire [7:0] _T_24780;
  wire [7:0] _T_24782;
  wire [7:0] _T_24784;
  wire [7:0] _T_24786;
  wire [7:0] _T_24788;
  wire [7:0] _T_24790;
  wire [7:0] _T_24792;
  wire [7:0] _T_24794;
  wire [7:0] _T_24796;
  wire [7:0] _T_24798;
  wire [7:0] _T_24800;
  wire [7:0] _T_24802;
  wire [7:0] _T_24804;
  wire [7:0] _T_24806;
  wire [7:0] _T_24808;
  wire [7:0] _T_24810;
  wire [7:0] _T_24812;
  wire [7:0] _T_24814;
  wire [7:0] _T_24816;
  wire [7:0] _T_24818;
  wire [7:0] _T_24820;
  wire [7:0] _T_24822;
  wire [7:0] _T_24824;
  wire [7:0] _T_24826;
  wire [7:0] _T_24828;
  wire [7:0] _T_24830;
  wire [7:0] _T_24832;
  wire [7:0] _T_24834;
  wire [7:0] _T_24836;
  wire [7:0] _T_24838;
  wire [7:0] _T_24840;
  wire [7:0] _T_24842;
  wire [7:0] _T_24844;
  wire [7:0] _T_24846;
  wire [7:0] _T_24848;
  wire [7:0] _T_24850;
  wire [7:0] _T_24852;
  wire [7:0] _T_24854;
  wire [7:0] _T_24856;
  wire [7:0] _T_24858;
  wire [7:0] _T_24860;
  wire [7:0] _T_24862;
  wire [7:0] _T_24864;
  wire [7:0] _T_24866;
  wire [7:0] _T_24868;
  wire [7:0] _T_24870;
  wire [7:0] _T_24872;
  wire [7:0] _T_24874;
  wire [7:0] _T_24876;
  wire [7:0] _T_24878;
  wire [7:0] _T_24880;
  wire [7:0] _T_24882;
  wire [7:0] _T_24884;
  wire [7:0] _T_24886;
  wire [7:0] _T_24888;
  wire [7:0] _T_24890;
  wire [7:0] _T_24892;
  wire [7:0] _T_24894;
  wire [7:0] _T_24896;
  wire [7:0] _T_24898;
  wire [7:0] _T_24900;
  wire [7:0] _T_24902;
  wire [7:0] _T_24904;
  wire [7:0] _T_24906;
  wire [7:0] _T_24908;
  wire [7:0] _T_24910;
  wire [7:0] _T_24912;
  wire [7:0] _T_24914;
  wire [7:0] _T_24916;
  wire [7:0] _T_24918;
  wire [7:0] _T_24920;
  wire [7:0] _T_24922;
  wire [7:0] _T_24924;
  wire [7:0] _T_24926;
  wire [7:0] _T_24928;
  wire [7:0] _T_24930;
  wire [7:0] _T_24932;
  wire [7:0] _T_24934;
  wire [7:0] _T_24936;
  wire [7:0] _T_24938;
  wire [7:0] _T_24940;
  wire [7:0] _T_24942;
  wire [7:0] _T_24944;
  wire [7:0] _T_24946;
  wire [7:0] _T_24948;
  wire [7:0] _T_24950;
  wire [7:0] _T_24952;
  wire [7:0] _T_24954;
  wire [7:0] _T_24956;
  wire [7:0] _T_24958;
  wire [7:0] _T_24960;
  wire [7:0] _T_24962;
  wire [7:0] _T_24964;
  wire [7:0] _T_24966;
  wire [7:0] _T_24968;
  wire [7:0] _T_24970;
  wire [7:0] _T_24972;
  wire [7:0] _T_24974;
  wire [7:0] _T_24976;
  wire [7:0] _T_24978;
  wire [7:0] _T_24980;
  wire [7:0] _T_24982;
  wire [7:0] _T_24984;
  wire [7:0] _T_24986;
  wire [7:0] _T_24988;
  wire [7:0] _T_24990;
  wire [7:0] _T_24992;
  wire [7:0] _T_24994;
  wire [7:0] _T_24996;
  wire [7:0] _T_24998;
  wire [7:0] _T_25000;
  wire [7:0] _T_25002;
  wire [7:0] _T_25004;
  wire [7:0] _T_25006;
  wire [7:0] _T_25008;
  wire [7:0] _T_25010;
  wire [7:0] _T_25012;
  wire [7:0] _T_25014;
  wire [7:0] _T_25016;
  wire [7:0] _T_25018;
  wire [7:0] _T_25020;
  wire [7:0] _T_25022;
  wire [7:0] _T_25024;
  wire [7:0] _T_25026;
  wire [7:0] _T_25028;
  wire [7:0] _T_25030;
  wire [7:0] _T_25032;
  wire [7:0] _T_25034;
  wire [7:0] _T_25036;
  wire [7:0] _T_25038;
  wire [7:0] _T_25040;
  wire [7:0] _T_25042;
  wire [7:0] _T_25044;
  wire [7:0] _T_25046;
  wire [7:0] _T_25048;
  wire [7:0] _T_25050;
  wire [7:0] _T_25052;
  wire [7:0] _T_25054;
  wire [7:0] _T_25056;
  wire [7:0] _T_25058;
  wire [7:0] _T_25060;
  wire [7:0] _T_25062;
  wire [7:0] _T_25064;
  wire [7:0] _T_25066;
  wire [7:0] _T_25068;
  wire [7:0] _T_25070;
  wire [7:0] _T_25072;
  wire [7:0] _T_25074;
  wire [7:0] _T_25076;
  wire [7:0] _T_25078;
  wire [7:0] _T_25080;
  wire [7:0] _T_25082;
  wire [7:0] _T_25084;
  wire [7:0] _T_25086;
  wire [7:0] _T_25088;
  wire [7:0] _T_25090;
  wire [7:0] _T_25092;
  wire [7:0] _T_25094;
  wire [7:0] _T_25096;
  wire [7:0] _T_25098;
  wire [7:0] _T_25100;
  wire [7:0] _T_25102;
  wire [7:0] _T_25104;
  wire [7:0] _T_25106;
  wire [7:0] _T_25108;
  wire [7:0] _T_25110;
  wire [7:0] _T_25112;
  wire [7:0] _T_25114;
  wire [7:0] _T_25116;
  wire [7:0] _T_25118;
  wire [7:0] _T_25120;
  wire [7:0] _T_25122;
  wire [7:0] _T_25124;
  wire [7:0] _T_25126;
  wire [7:0] _T_25128;
  wire [7:0] _T_25130;
  wire [7:0] _T_25132;
  wire [7:0] _T_25134;
  wire [7:0] _T_25136;
  wire [7:0] _T_25138;
  wire [7:0] _T_25140;
  wire [7:0] _T_25142;
  wire [7:0] _T_25144;
  wire [7:0] _T_25146;
  wire [7:0] _T_25148;
  wire [7:0] _T_25150;
  wire [7:0] _T_25152;
  wire [7:0] _T_25154;
  wire [7:0] _T_25156;
  wire [7:0] _T_25158;
  wire [7:0] _T_25160;
  wire [7:0] _T_25162;
  wire [7:0] _T_25164;
  wire [7:0] _T_25166;
  wire [7:0] _T_25168;
  wire [7:0] _T_25170;
  wire [7:0] _T_25172;
  wire [7:0] _T_25174;
  wire [7:0] _T_25176;
  wire [7:0] _T_25178;
  wire [7:0] _T_25180;
  wire [7:0] _T_25182;
  wire [7:0] _T_25184;
  wire [7:0] _T_25186;
  wire [7:0] _T_25188;
  wire [7:0] _T_25190;
  wire [7:0] _T_25192;
  wire [7:0] _T_25194;
  wire [7:0] _T_25196;
  wire [7:0] _T_25198;
  wire [7:0] _T_25200;
  wire [7:0] _T_25202;
  wire [7:0] _T_25204;
  wire [7:0] _T_25206;
  wire [7:0] _T_25208;
  wire [7:0] _T_25210;
  wire [7:0] _T_25212;
  wire [7:0] _T_25214;
  wire [7:0] _T_25216;
  wire [7:0] _T_25218;
  wire [7:0] _T_25220;
  wire [7:0] _T_25222;
  wire [7:0] _T_25224;
  wire [7:0] _T_25226;
  wire [7:0] _T_25228;
  wire [7:0] _T_25230;
  wire [7:0] _T_25232;
  wire [7:0] _T_25234;
  wire [7:0] _T_25236;
  wire [7:0] _T_25238;
  wire [7:0] _T_25240;
  wire [7:0] _T_25242;
  wire [7:0] _T_25244;
  wire [7:0] _T_25246;
  wire [7:0] _T_25248;
  wire [7:0] _T_25250;
  wire [7:0] _T_25252;
  wire [7:0] _T_25254;
  wire [7:0] _T_25256;
  wire [7:0] _T_25258;
  wire [7:0] _T_25260;
  wire [7:0] _T_25262;
  wire [7:0] _T_25264;
  wire [7:0] _T_25266;
  wire [7:0] _T_25268;
  wire [7:0] _T_25270;
  wire [7:0] _T_25272;
  wire [7:0] _T_25274;
  wire [7:0] _T_25276;
  wire [7:0] _T_25278;
  wire [7:0] _T_25280;
  wire [7:0] _T_25282;
  wire [7:0] _T_25284;
  wire [7:0] _T_25286;
  wire [7:0] _T_25288;
  wire [7:0] _T_25290;
  wire [7:0] _T_25292;
  wire [7:0] _T_25294;
  wire [7:0] _T_25296;
  wire [7:0] _T_25298;
  wire [7:0] _T_25300;
  wire [7:0] _T_25302;
  wire [7:0] _T_25304;
  wire [7:0] _T_25306;
  wire [7:0] _T_25308;
  wire [7:0] _T_25310;
  wire [7:0] _T_25312;
  wire [7:0] _T_25314;
  wire [7:0] _T_25316;
  wire [7:0] _T_25318;
  wire [7:0] _T_25320;
  wire [7:0] _T_25322;
  wire [7:0] _T_25324;
  wire [7:0] _T_25326;
  wire [7:0] _T_25328;
  wire [7:0] _T_25330;
  wire [7:0] _T_25332;
  wire [7:0] _T_25334;
  wire [7:0] _T_25336;
  wire [7:0] _T_25338;
  wire [7:0] _T_25340;
  wire [7:0] _T_25342;
  wire [7:0] _T_25344;
  wire [7:0] _T_25346;
  wire [7:0] _T_25348;
  wire [7:0] _T_25350;
  wire [7:0] _T_25352;
  wire [7:0] _T_25354;
  wire [7:0] _T_25356;
  wire [7:0] _T_25358;
  wire [7:0] _T_25360;
  wire [7:0] _T_25362;
  wire [7:0] _T_25364;
  wire [7:0] _T_25366;
  wire [7:0] _T_25368;
  wire [7:0] _T_25370;
  wire [7:0] _T_25372;
  wire [7:0] _T_25374;
  wire [7:0] _T_25376;
  wire [7:0] _T_25378;
  wire [7:0] _T_25380;
  wire [7:0] _T_25382;
  wire [7:0] _T_25384;
  wire [7:0] _T_25386;
  wire [7:0] _T_25388;
  wire [7:0] _T_25390;
  wire [7:0] _T_25392;
  wire [7:0] _T_25394;
  wire [7:0] _T_25396;
  wire [7:0] _T_25398;
  wire [7:0] _T_25400;
  wire [7:0] _T_25402;
  wire [7:0] _T_25404;
  wire [7:0] _T_25406;
  wire [7:0] _T_25408;
  wire [7:0] _T_25410;
  wire [7:0] _T_25412;
  wire [7:0] _T_25414;
  wire [7:0] _T_25416;
  wire [7:0] _T_25418;
  wire [7:0] _T_25420;
  wire [7:0] _T_25422;
  wire [7:0] _T_25424;
  wire [7:0] _T_25426;
  wire [7:0] _T_25428;
  wire [7:0] _T_25430;
  wire [7:0] _T_25432;
  wire [7:0] _T_25434;
  wire [7:0] _T_25436;
  wire [7:0] _T_25438;
  wire [7:0] _T_25440;
  wire [7:0] _T_25442;
  wire [7:0] _T_25444;
  wire [7:0] _T_25446;
  wire [7:0] _T_25448;
  wire [7:0] _T_25450;
  wire [7:0] _T_25452;
  wire [7:0] _T_25454;
  wire [7:0] _T_25456;
  wire [7:0] _T_25458;
  wire [7:0] _T_25460;
  wire [7:0] _T_25462;
  wire [7:0] _T_25464;
  wire [7:0] _T_25466;
  wire [7:0] _T_25468;
  wire [7:0] _T_25470;
  wire [7:0] _T_25472;
  wire [7:0] _T_25474;
  wire [7:0] _T_25476;
  wire [7:0] _T_25478;
  wire [7:0] _T_25480;
  wire [7:0] _T_25482;
  wire [7:0] _T_25484;
  wire [7:0] _T_25486;
  wire [7:0] _T_25488;
  wire [7:0] _T_25490;
  wire [7:0] _T_25492;
  wire [7:0] _T_25494;
  wire [7:0] _T_25496;
  wire [7:0] _T_25498;
  wire [7:0] _T_25500;
  wire [7:0] _T_25502;
  wire [7:0] _T_25504;
  wire [7:0] _T_25506;
  wire [7:0] _T_25508;
  wire [7:0] _T_25510;
  wire [7:0] _T_25512;
  wire [7:0] _T_25514;
  wire [7:0] _T_25516;
  wire [7:0] _T_25518;
  wire [7:0] _T_25520;
  wire [7:0] _T_25522;
  wire [7:0] _T_25524;
  wire [7:0] _T_25526;
  wire [7:0] _T_25528;
  wire [7:0] _T_25530;
  wire [7:0] _T_25532;
  wire [7:0] _T_25534;
  wire [7:0] _T_25536;
  wire [7:0] _T_25538;
  wire [7:0] _T_25540;
  wire [7:0] _T_25542;
  wire [7:0] _T_25544;
  wire [7:0] _T_25546;
  wire [7:0] _T_25548;
  wire [7:0] _T_25550;
  wire [7:0] _T_25552;
  wire [7:0] _T_25554;
  wire [7:0] _T_25556;
  wire [7:0] _T_25558;
  wire [7:0] _T_25560;
  wire [7:0] _T_25562;
  wire [7:0] _T_25564;
  wire [7:0] _T_25566;
  wire [7:0] _T_25568;
  wire [7:0] _T_25570;
  wire [7:0] _T_25572;
  wire [7:0] _T_25574;
  wire [7:0] _T_25576;
  wire [7:0] _T_25578;
  wire [7:0] _T_25580;
  wire [7:0] _T_25582;
  wire [7:0] _T_25584;
  wire [7:0] _T_25586;
  wire [7:0] _T_25588;
  wire [7:0] _T_25590;
  wire [7:0] _T_25592;
  wire [7:0] _T_25594;
  wire [7:0] _T_25596;
  wire [7:0] _T_25598;
  wire [7:0] _T_25600;
  wire [7:0] _T_25602;
  wire [7:0] _T_25604;
  wire [7:0] _T_25606;
  wire [7:0] _T_25608;
  wire [7:0] _T_25610;
  wire [7:0] _T_25612;
  wire [7:0] _T_25614;
  wire [7:0] _T_25616;
  wire [7:0] _T_25618;
  wire [7:0] _T_25620;
  wire [7:0] _T_25622;
  wire [7:0] _T_25624;
  wire [7:0] _T_25626;
  wire [7:0] _T_25628;
  wire [7:0] _T_25630;
  wire [7:0] _T_25632;
  wire [7:0] _T_25634;
  wire [7:0] _T_25636;
  wire [7:0] _T_25638;
  wire [7:0] _T_25640;
  wire [7:0] _T_25642;
  wire [7:0] _T_25644;
  wire [7:0] _T_25646;
  wire [7:0] _T_25648;
  wire [7:0] _T_25650;
  wire [7:0] _T_25652;
  wire [7:0] _T_25654;
  wire [7:0] _T_25656;
  wire [7:0] _T_25658;
  wire [7:0] _T_25660;
  wire [7:0] _T_25662;
  wire [7:0] _T_25664;
  wire [7:0] _T_25666;
  wire [7:0] _T_25668;
  wire [7:0] _T_25670;
  wire [7:0] _T_25672;
  wire [7:0] _T_25674;
  wire [7:0] _T_25676;
  wire [7:0] _T_25678;
  wire [7:0] _T_25680;
  wire [7:0] _T_25682;
  wire [7:0] _T_25684;
  wire [7:0] _T_25686;
  wire [7:0] _T_25688;
  wire [7:0] _T_25690;
  wire [7:0] _T_25692;
  wire [7:0] _T_25694;
  wire [7:0] _T_25696;
  wire [7:0] _T_25698;
  wire [7:0] _T_25700;
  wire [7:0] _T_25702;
  wire [7:0] _T_25704;
  wire [7:0] _T_25706;
  wire [7:0] _T_25708;
  wire [7:0] _T_25710;
  wire [7:0] _T_25712;
  wire [7:0] _T_25714;
  wire [7:0] _T_25716;
  wire [7:0] _T_25718;
  wire [7:0] _T_25720;
  wire [7:0] _T_25722;
  wire [7:0] _T_25724;
  wire [7:0] _T_25726;
  wire [7:0] _T_25728;
  wire [7:0] _T_25730;
  wire [7:0] _T_25732;
  wire [7:0] _T_25734;
  wire [7:0] _T_25736;
  wire [7:0] _T_25738;
  wire [7:0] _T_25740;
  wire [7:0] _T_25742;
  wire [7:0] _T_25744;
  wire [7:0] _T_25746;
  wire [7:0] _T_25748;
  wire [7:0] _T_25750;
  wire [7:0] _T_25752;
  wire [7:0] _T_25754;
  wire [7:0] _T_25756;
  wire [7:0] _T_25758;
  wire [7:0] _T_25760;
  wire [7:0] _T_25762;
  wire [7:0] _T_25764;
  wire [7:0] _T_25766;
  wire [7:0] _T_25768;
  wire [7:0] _T_25770;
  wire [7:0] _T_25772;
  wire [7:0] _T_25774;
  wire [7:0] _T_25776;
  wire [7:0] _T_25778;
  wire [7:0] _T_25780;
  wire [7:0] _T_25782;
  wire [7:0] _T_25784;
  wire [7:0] _T_25786;
  wire [7:0] _T_25788;
  wire [7:0] _T_25790;
  wire [7:0] _T_25792;
  wire  _T_25899;
  wire [9:0] _T_25900;
  wire [11:0] _T_25901;
  wire [9:0] _T_26947;
  wire [9:0] _T_26948;
  wire  _T_26950;
  wire [9:0] _T_26956;
  wire [9:0] _T_26957;
  wire  _T_26959;
  wire [9:0] _T_26965;
  wire [9:0] _T_26966;
  wire  _T_26968;
  wire [9:0] _T_26974;
  wire [9:0] _T_26975;
  wire  _T_26977;
  wire [9:0] _T_26983;
  wire [9:0] _T_26984;
  wire  _T_26986;
  wire [9:0] _T_26992;
  wire [9:0] _T_26993;
  wire  _T_26995;
  wire [9:0] _T_27001;
  wire [9:0] _T_27002;
  wire  _T_27004;
  wire [9:0] _T_27010;
  wire [9:0] _T_27011;
  wire  _T_27013;
  wire [9:0] _T_27019;
  wire [9:0] _T_27020;
  wire  _T_27022;
  wire [9:0] _T_27028;
  wire [9:0] _T_27029;
  wire  _T_27031;
  wire [9:0] _T_27037;
  wire [9:0] _T_27038;
  wire  _T_27040;
  wire [9:0] _T_27046;
  wire [9:0] _T_27047;
  wire  _T_27049;
  wire [9:0] _T_27055;
  wire [9:0] _T_27056;
  wire  _T_27058;
  wire [9:0] _T_27064;
  wire [9:0] _T_27065;
  wire  _T_27067;
  wire [9:0] _T_27073;
  wire [9:0] _T_27074;
  wire  _T_27076;
  wire [9:0] _T_27082;
  wire [9:0] _T_27083;
  wire  _T_27085;
  wire [9:0] _T_27091;
  wire [9:0] _T_27092;
  wire  _T_27094;
  wire [9:0] _T_27100;
  wire [9:0] _T_27101;
  wire  _T_27103;
  wire [9:0] _T_27109;
  wire [9:0] _T_27110;
  wire  _T_27112;
  wire [9:0] _T_27118;
  wire [9:0] _T_27119;
  wire  _T_27121;
  wire [9:0] _T_27127;
  wire [9:0] _T_27128;
  wire  _T_27130;
  wire [9:0] _T_27136;
  wire [9:0] _T_27137;
  wire  _T_27139;
  wire [9:0] _T_27145;
  wire [9:0] _T_27146;
  wire  _T_27148;
  wire [9:0] _T_27154;
  wire [9:0] _T_27155;
  wire  _T_27157;
  wire [9:0] _T_27163;
  wire [9:0] _T_27164;
  wire  _T_27166;
  wire [9:0] _T_27172;
  wire [9:0] _T_27173;
  wire  _T_27175;
  wire [9:0] _T_27181;
  wire [9:0] _T_27182;
  wire  _T_27184;
  wire [9:0] _T_27190;
  wire [9:0] _T_27191;
  wire  _T_27193;
  wire [9:0] _T_27199;
  wire [9:0] _T_27200;
  wire  _T_27202;
  wire [9:0] _T_27208;
  wire [9:0] _T_27209;
  wire  _T_27211;
  wire [9:0] _T_27217;
  wire [9:0] _T_27218;
  wire  _T_27220;
  wire [9:0] _T_27226;
  wire [9:0] _T_27227;
  wire  _T_27229;
  wire [9:0] _T_27235;
  wire [9:0] _T_27236;
  wire  _T_27238;
  wire [9:0] _T_27244;
  wire [9:0] _T_27245;
  wire  _T_27247;
  wire [9:0] _T_27253;
  wire [9:0] _T_27254;
  wire  _T_27256;
  wire [9:0] _T_27262;
  wire [9:0] _T_27263;
  wire  _T_27265;
  wire [9:0] _T_27271;
  wire [9:0] _T_27272;
  wire  _T_27274;
  wire [9:0] _T_27280;
  wire [9:0] _T_27281;
  wire  _T_27283;
  wire [9:0] _T_27289;
  wire [9:0] _T_27290;
  wire  _T_27292;
  wire [9:0] _T_27298;
  wire [9:0] _T_27299;
  wire  _T_27301;
  wire [9:0] _T_27307;
  wire [9:0] _T_27308;
  wire  _T_27310;
  wire [9:0] _T_27316;
  wire [9:0] _T_27317;
  wire  _T_27319;
  wire [9:0] _T_27325;
  wire [9:0] _T_27326;
  wire  _T_27328;
  wire [9:0] _T_27334;
  wire [9:0] _T_27335;
  wire  _T_27337;
  wire [9:0] _T_27343;
  wire [9:0] _T_27344;
  wire  _T_27346;
  wire [9:0] _T_27352;
  wire [9:0] _T_27353;
  wire  _T_27355;
  wire [9:0] _T_27361;
  wire [9:0] _T_27362;
  wire  _T_27364;
  wire [9:0] _T_27370;
  wire [9:0] _T_27371;
  wire  _T_27373;
  wire [9:0] _T_27379;
  wire [9:0] _T_27380;
  wire  _T_27382;
  wire [9:0] _T_27388;
  wire [9:0] _T_27389;
  wire  _T_27391;
  wire [9:0] _T_27397;
  wire [9:0] _T_27398;
  wire  _T_27400;
  wire [9:0] _T_27406;
  wire [9:0] _T_27407;
  wire  _T_27409;
  wire [9:0] _T_27415;
  wire [9:0] _T_27416;
  wire  _T_27418;
  wire [9:0] _T_27424;
  wire [9:0] _T_27425;
  wire  _T_27427;
  wire [9:0] _T_27433;
  wire [9:0] _T_27434;
  wire  _T_27436;
  wire [9:0] _T_27442;
  wire [9:0] _T_27443;
  wire  _T_27445;
  wire [9:0] _T_27451;
  wire [9:0] _T_27452;
  wire  _T_27454;
  wire [9:0] _T_27460;
  wire [9:0] _T_27461;
  wire  _T_27463;
  wire [9:0] _T_27469;
  wire [9:0] _T_27470;
  wire  _T_27472;
  wire [9:0] _T_27478;
  wire [9:0] _T_27479;
  wire  _T_27481;
  wire [9:0] _T_27487;
  wire [9:0] _T_27488;
  wire  _T_27490;
  wire [9:0] _T_27496;
  wire [9:0] _T_27497;
  wire  _T_27499;
  wire [9:0] _T_27505;
  wire [9:0] _T_27506;
  wire  _T_27508;
  wire [9:0] _T_27514;
  wire [9:0] _T_27515;
  wire  _T_27517;
  wire [9:0] _T_27523;
  wire [9:0] _T_27524;
  wire  _T_27526;
  wire [9:0] _T_27532;
  wire [9:0] _T_27533;
  wire  _T_27535;
  wire [9:0] _T_27541;
  wire [9:0] _T_27542;
  wire  _T_27544;
  wire [9:0] _T_27550;
  wire [9:0] _T_27551;
  wire  _T_27553;
  wire [9:0] _T_27559;
  wire [9:0] _T_27560;
  wire  _T_27562;
  wire [9:0] _T_27568;
  wire [9:0] _T_27569;
  wire  _T_27571;
  wire [9:0] _T_27577;
  wire [9:0] _T_27578;
  wire  _T_27580;
  wire [9:0] _T_27586;
  wire [9:0] _T_27587;
  wire  _T_27589;
  wire [9:0] _T_27595;
  wire [9:0] _T_27596;
  wire  _T_27598;
  wire [9:0] _T_27604;
  wire [9:0] _T_27605;
  wire  _T_27607;
  wire [9:0] _T_27613;
  wire [9:0] _T_27614;
  wire  _T_27616;
  wire [9:0] _T_27622;
  wire [9:0] _T_27623;
  wire  _T_27625;
  wire [9:0] _T_27631;
  wire [9:0] _T_27632;
  wire  _T_27634;
  wire [9:0] _T_27640;
  wire [9:0] _T_27641;
  wire  _T_27643;
  wire [9:0] _T_27649;
  wire [9:0] _T_27650;
  wire  _T_27652;
  wire [9:0] _T_27658;
  wire [9:0] _T_27659;
  wire  _T_27661;
  wire [9:0] _T_27667;
  wire [9:0] _T_27668;
  wire  _T_27670;
  wire [9:0] _T_27676;
  wire [9:0] _T_27677;
  wire  _T_27679;
  wire [9:0] _T_27685;
  wire [9:0] _T_27686;
  wire  _T_27688;
  wire [9:0] _T_27694;
  wire [9:0] _T_27695;
  wire  _T_27697;
  wire [9:0] _T_27703;
  wire [9:0] _T_27704;
  wire  _T_27706;
  wire [9:0] _T_27712;
  wire [9:0] _T_27713;
  wire  _T_27715;
  wire [9:0] _T_27721;
  wire [9:0] _T_27722;
  wire  _T_27724;
  wire [9:0] _T_27730;
  wire [9:0] _T_27731;
  wire  _T_27733;
  wire [9:0] _T_27739;
  wire [9:0] _T_27740;
  wire  _T_27742;
  wire [9:0] _T_27748;
  wire [9:0] _T_27749;
  wire  _T_27751;
  wire [9:0] _T_27757;
  wire [9:0] _T_27758;
  wire  _T_27760;
  wire [9:0] _T_27766;
  wire [9:0] _T_27767;
  wire  _T_27769;
  wire [9:0] _T_27775;
  wire [9:0] _T_27776;
  wire  _T_27778;
  wire [9:0] _T_27784;
  wire [9:0] _T_27785;
  wire  _T_27787;
  wire [9:0] _T_27793;
  wire [9:0] _T_27794;
  wire  _T_27796;
  wire [9:0] _T_27802;
  wire [9:0] _T_27803;
  wire  _T_27805;
  wire [9:0] _T_27811;
  wire [9:0] _T_27812;
  wire  _T_27814;
  wire [9:0] _T_27820;
  wire [9:0] _T_27821;
  wire  _T_27823;
  wire [9:0] _T_27829;
  wire [9:0] _T_27830;
  wire  _T_27832;
  wire [9:0] _T_27838;
  wire [9:0] _T_27839;
  wire  _T_27841;
  wire [9:0] _T_27847;
  wire [9:0] _T_27848;
  wire  _T_27850;
  wire [9:0] _T_27856;
  wire [9:0] _T_27857;
  wire  _T_27859;
  wire [9:0] _T_27865;
  wire [9:0] _T_27866;
  wire  _T_27868;
  wire [9:0] _T_27874;
  wire [9:0] _T_27875;
  wire  _T_27877;
  wire [9:0] _T_27883;
  wire [9:0] _T_27884;
  wire  _T_27886;
  wire [9:0] _T_27892;
  wire [9:0] _T_27893;
  wire  _T_27895;
  wire [9:0] _T_27901;
  wire [9:0] _T_27902;
  wire  _T_27904;
  wire [9:0] _T_27910;
  wire [9:0] _T_27911;
  wire  _T_27913;
  wire [9:0] _T_27919;
  wire [9:0] _T_27920;
  wire  _T_27922;
  wire [9:0] _T_27928;
  wire [9:0] _T_27929;
  wire  _T_27931;
  wire [9:0] _T_27937;
  wire [9:0] _T_27938;
  wire  _T_27940;
  wire [9:0] _T_27946;
  wire [9:0] _T_27947;
  wire  _T_27949;
  wire [9:0] _T_27955;
  wire [9:0] _T_27956;
  wire  _T_27958;
  wire [9:0] _T_27964;
  wire [9:0] _T_27965;
  wire  _T_27967;
  wire [9:0] _T_27973;
  wire [9:0] _T_27974;
  wire  _T_27976;
  wire [9:0] _T_27982;
  wire [9:0] _T_27983;
  wire  _T_27985;
  wire [9:0] _T_27991;
  wire [9:0] _T_27992;
  wire  _T_27994;
  wire [9:0] _T_28000;
  wire [9:0] _T_28001;
  wire  _T_28003;
  wire [9:0] _T_28009;
  wire [9:0] _T_28010;
  wire  _T_28012;
  wire [9:0] _T_28018;
  wire [9:0] _T_28019;
  wire  _T_28021;
  wire [9:0] _T_28027;
  wire [9:0] _T_28028;
  wire  _T_28030;
  wire [9:0] _T_28036;
  wire [9:0] _T_28037;
  wire  _T_28039;
  wire [9:0] _T_28045;
  wire [9:0] _T_28046;
  wire  _T_28048;
  wire [9:0] _T_28054;
  wire [9:0] _T_28055;
  wire  _T_28057;
  wire [9:0] _T_28063;
  wire [9:0] _T_28064;
  wire  _T_28066;
  wire [9:0] _T_28072;
  wire [9:0] _T_28073;
  wire  _T_28075;
  wire [9:0] _T_28081;
  wire [9:0] _T_28082;
  wire  _T_28084;
  wire [9:0] _T_28090;
  wire [9:0] _T_28091;
  wire  _T_28093;
  wire [9:0] _T_28099;
  wire [9:0] _T_28100;
  wire  _T_28102;
  wire [9:0] _T_28108;
  wire [9:0] _T_28109;
  wire  _T_28111;
  wire [9:0] _T_28117;
  wire [9:0] _T_28118;
  wire  _T_28120;
  wire [9:0] _T_28126;
  wire [9:0] _T_28127;
  wire  _T_28129;
  wire [9:0] _T_28135;
  wire [9:0] _T_28136;
  wire  _T_28138;
  wire [9:0] _T_28144;
  wire [9:0] _T_28145;
  wire  _T_28147;
  wire [9:0] _T_28153;
  wire [9:0] _T_28154;
  wire  _T_28156;
  wire [9:0] _T_28162;
  wire [9:0] _T_28163;
  wire  _T_28165;
  wire [9:0] _T_28171;
  wire [9:0] _T_28172;
  wire  _T_28174;
  wire [9:0] _T_28180;
  wire [9:0] _T_28181;
  wire  _T_28183;
  wire [9:0] _T_28189;
  wire [9:0] _T_28190;
  wire  _T_28192;
  wire [9:0] _T_28198;
  wire [9:0] _T_28199;
  wire  _T_28201;
  wire [9:0] _T_28207;
  wire [9:0] _T_28208;
  wire  _T_28210;
  wire [9:0] _T_28216;
  wire [9:0] _T_28217;
  wire  _T_28219;
  wire [9:0] _T_28225;
  wire [9:0] _T_28226;
  wire  _T_28228;
  wire [9:0] _T_28234;
  wire [9:0] _T_28235;
  wire  _T_28237;
  wire [9:0] _T_28243;
  wire [9:0] _T_28244;
  wire  _T_28246;
  wire [9:0] _T_28252;
  wire [9:0] _T_28253;
  wire  _T_28255;
  wire [9:0] _T_28261;
  wire [9:0] _T_28262;
  wire  _T_28264;
  wire [9:0] _T_28270;
  wire [9:0] _T_28271;
  wire  _T_28273;
  wire [9:0] _T_28279;
  wire [9:0] _T_28280;
  wire  _T_28282;
  wire [9:0] _T_28288;
  wire [9:0] _T_28289;
  wire  _T_28291;
  wire [9:0] _T_28297;
  wire [9:0] _T_28298;
  wire  _T_28300;
  wire [9:0] _T_28306;
  wire [9:0] _T_28307;
  wire  _T_28309;
  wire [9:0] _T_28315;
  wire [9:0] _T_28316;
  wire  _T_28318;
  wire [9:0] _T_28324;
  wire [9:0] _T_28325;
  wire  _T_28327;
  wire [9:0] _T_28333;
  wire [9:0] _T_28334;
  wire  _T_28336;
  wire [9:0] _T_28342;
  wire [9:0] _T_28343;
  wire  _T_28345;
  wire [9:0] _T_28351;
  wire [9:0] _T_28352;
  wire  _T_28354;
  wire [9:0] _T_28360;
  wire [9:0] _T_28361;
  wire  _T_28363;
  wire [9:0] _T_28369;
  wire [9:0] _T_28370;
  wire  _T_28372;
  wire [9:0] _T_28378;
  wire [9:0] _T_28379;
  wire  _T_28381;
  wire [9:0] _T_28387;
  wire [9:0] _T_28388;
  wire  _T_28390;
  wire [9:0] _T_28396;
  wire [9:0] _T_28397;
  wire  _T_28399;
  wire [9:0] _T_28405;
  wire [9:0] _T_28406;
  wire  _T_28408;
  wire [9:0] _T_28414;
  wire [9:0] _T_28415;
  wire  _T_28417;
  wire [9:0] _T_28423;
  wire [9:0] _T_28424;
  wire  _T_28426;
  wire [9:0] _T_28432;
  wire [9:0] _T_28433;
  wire  _T_28435;
  wire [9:0] _T_28441;
  wire [9:0] _T_28442;
  wire  _T_28444;
  wire [9:0] _T_28450;
  wire [9:0] _T_28451;
  wire  _T_28453;
  wire [9:0] _T_28459;
  wire [9:0] _T_28460;
  wire  _T_28462;
  wire [9:0] _T_28468;
  wire [9:0] _T_28469;
  wire  _T_28471;
  wire [9:0] _T_28477;
  wire [9:0] _T_28478;
  wire  _T_28480;
  wire [9:0] _T_28486;
  wire [9:0] _T_28487;
  wire  _T_28489;
  wire [9:0] _T_28495;
  wire [9:0] _T_28496;
  wire  _T_28498;
  wire [9:0] _T_28504;
  wire [9:0] _T_28505;
  wire  _T_28507;
  wire [9:0] _T_28513;
  wire [9:0] _T_28514;
  wire  _T_28516;
  wire [9:0] _T_28522;
  wire [9:0] _T_28523;
  wire  _T_28525;
  wire [9:0] _T_28531;
  wire [9:0] _T_28532;
  wire  _T_28534;
  wire [9:0] _T_28540;
  wire [9:0] _T_28541;
  wire  _T_28543;
  wire [9:0] _T_28549;
  wire [9:0] _T_28550;
  wire  _T_28552;
  wire [9:0] _T_28558;
  wire [9:0] _T_28559;
  wire  _T_28561;
  wire [9:0] _T_28567;
  wire [9:0] _T_28568;
  wire  _T_28570;
  wire [9:0] _T_28576;
  wire [9:0] _T_28577;
  wire  _T_28579;
  wire [9:0] _T_28585;
  wire [9:0] _T_28586;
  wire  _T_28588;
  wire [9:0] _T_28594;
  wire [9:0] _T_28595;
  wire  _T_28597;
  wire [9:0] _T_28603;
  wire [9:0] _T_28604;
  wire  _T_28606;
  wire [9:0] _T_28612;
  wire [9:0] _T_28613;
  wire  _T_28615;
  wire [9:0] _T_28621;
  wire [9:0] _T_28622;
  wire  _T_28624;
  wire [9:0] _T_28630;
  wire [9:0] _T_28631;
  wire  _T_28633;
  wire [9:0] _T_28639;
  wire [9:0] _T_28640;
  wire  _T_28642;
  wire [9:0] _T_28648;
  wire [9:0] _T_28649;
  wire  _T_28651;
  wire [9:0] _T_28657;
  wire [9:0] _T_28658;
  wire  _T_28660;
  wire [9:0] _T_28666;
  wire [9:0] _T_28667;
  wire  _T_28669;
  wire [9:0] _T_28675;
  wire [9:0] _T_28676;
  wire  _T_28678;
  wire [9:0] _T_28684;
  wire [9:0] _T_28685;
  wire  _T_28687;
  wire [9:0] _T_28693;
  wire [9:0] _T_28694;
  wire  _T_28696;
  wire [9:0] _T_28702;
  wire [9:0] _T_28703;
  wire  _T_28705;
  wire [9:0] _T_28711;
  wire [9:0] _T_28712;
  wire  _T_28714;
  wire [9:0] _T_28720;
  wire [9:0] _T_28721;
  wire  _T_28723;
  wire [9:0] _T_28729;
  wire [9:0] _T_28730;
  wire  _T_28732;
  wire [9:0] _T_28738;
  wire [9:0] _T_28739;
  wire  _T_28741;
  wire [9:0] _T_28747;
  wire [9:0] _T_28748;
  wire  _T_28750;
  wire [9:0] _T_28756;
  wire [9:0] _T_28757;
  wire  _T_28759;
  wire [9:0] _T_28765;
  wire [9:0] _T_28766;
  wire  _T_28768;
  wire [9:0] _T_28774;
  wire [9:0] _T_28775;
  wire  _T_28777;
  wire [9:0] _T_28783;
  wire [9:0] _T_28784;
  wire  _T_28786;
  wire [9:0] _T_28792;
  wire [9:0] _T_28793;
  wire  _T_28795;
  wire [9:0] _T_28801;
  wire [9:0] _T_28802;
  wire  _T_28804;
  wire [9:0] _T_28810;
  wire [9:0] _T_28811;
  wire  _T_28813;
  wire [9:0] _T_28819;
  wire [9:0] _T_28820;
  wire  _T_28822;
  wire [9:0] _T_28828;
  wire [9:0] _T_28829;
  wire  _T_28831;
  wire [9:0] _T_28837;
  wire [9:0] _T_28838;
  wire  _T_28840;
  wire [9:0] _T_28846;
  wire [9:0] _T_28847;
  wire  _T_28849;
  wire [9:0] _T_28855;
  wire [9:0] _T_28856;
  wire  _T_28858;
  wire [9:0] _T_28864;
  wire [9:0] _T_28865;
  wire  _T_28867;
  wire [9:0] _T_28873;
  wire [9:0] _T_28874;
  wire  _T_28876;
  wire [9:0] _T_28882;
  wire [9:0] _T_28883;
  wire  _T_28885;
  wire [9:0] _T_28891;
  wire [9:0] _T_28892;
  wire  _T_28894;
  wire [9:0] _T_28900;
  wire [9:0] _T_28901;
  wire  _T_28903;
  wire [9:0] _T_28909;
  wire [9:0] _T_28910;
  wire  _T_28912;
  wire [9:0] _T_28918;
  wire [9:0] _T_28919;
  wire  _T_28921;
  wire [9:0] _T_28927;
  wire [9:0] _T_28928;
  wire  _T_28930;
  wire [9:0] _T_28936;
  wire [9:0] _T_28937;
  wire  _T_28939;
  wire [9:0] _T_28945;
  wire [9:0] _T_28946;
  wire  _T_28948;
  wire [9:0] _T_28954;
  wire [9:0] _T_28955;
  wire  _T_28957;
  wire [9:0] _T_28963;
  wire [9:0] _T_28964;
  wire  _T_28966;
  wire [9:0] _T_28972;
  wire [9:0] _T_28973;
  wire  _T_28975;
  wire [9:0] _T_28981;
  wire [9:0] _T_28982;
  wire  _T_28984;
  wire [9:0] _T_28990;
  wire [9:0] _T_28991;
  wire  _T_28993;
  wire [9:0] _T_28999;
  wire [9:0] _T_29000;
  wire  _T_29002;
  wire [9:0] _T_29008;
  wire [9:0] _T_29009;
  wire  _T_29011;
  wire [9:0] _T_29017;
  wire [9:0] _T_29018;
  wire  _T_29020;
  wire [9:0] _T_29026;
  wire [9:0] _T_29027;
  wire  _T_29029;
  wire [9:0] _T_29035;
  wire [9:0] _T_29036;
  wire  _T_29038;
  wire [9:0] _T_29044;
  wire [9:0] _T_29045;
  wire  _T_29047;
  wire [9:0] _T_29053;
  wire [9:0] _T_29054;
  wire  _T_29056;
  wire [9:0] _T_29062;
  wire [9:0] _T_29063;
  wire  _T_29065;
  wire [9:0] _T_29071;
  wire [9:0] _T_29072;
  wire  _T_29074;
  wire [9:0] _T_29080;
  wire [9:0] _T_29081;
  wire  _T_29083;
  wire [9:0] _T_29089;
  wire [9:0] _T_29090;
  wire  _T_29092;
  wire [9:0] _T_29098;
  wire [9:0] _T_29099;
  wire  _T_29101;
  wire [9:0] _T_29107;
  wire [9:0] _T_29108;
  wire  _T_29110;
  wire [9:0] _T_29116;
  wire [9:0] _T_29117;
  wire  _T_29119;
  wire [9:0] _T_29125;
  wire [9:0] _T_29126;
  wire  _T_29128;
  wire [9:0] _T_29134;
  wire [9:0] _T_29135;
  wire  _T_29137;
  wire [9:0] _T_29143;
  wire [9:0] _T_29144;
  wire  _T_29146;
  wire [9:0] _T_29152;
  wire [9:0] _T_29153;
  wire  _T_29155;
  wire [9:0] _T_29161;
  wire [9:0] _T_29162;
  wire  _T_29164;
  wire [9:0] _T_29170;
  wire [9:0] _T_29171;
  wire  _T_29173;
  wire [9:0] _T_29179;
  wire [9:0] _T_29180;
  wire  _T_29182;
  wire [9:0] _T_29188;
  wire [9:0] _T_29189;
  wire  _T_29191;
  wire [9:0] _T_29197;
  wire [9:0] _T_29198;
  wire  _T_29200;
  wire [9:0] _T_29206;
  wire [9:0] _T_29207;
  wire  _T_29209;
  wire [9:0] _T_29215;
  wire [9:0] _T_29216;
  wire  _T_29218;
  wire [9:0] _T_29224;
  wire [9:0] _T_29225;
  wire  _T_29227;
  wire [9:0] _T_29233;
  wire [9:0] _T_29234;
  wire  _T_29236;
  wire [9:0] _T_29242;
  wire [9:0] _T_29243;
  wire  _T_29245;
  wire [9:0] _T_29251;
  wire [9:0] _T_29252;
  wire  _T_29254;
  wire [9:0] _T_29260;
  wire [9:0] _T_29261;
  wire  _T_29263;
  wire [9:0] _T_29269;
  wire [9:0] _T_29270;
  wire  _T_29272;
  wire [9:0] _T_29278;
  wire [9:0] _T_29279;
  wire  _T_29281;
  wire [9:0] _T_29287;
  wire [9:0] _T_29288;
  wire  _T_29290;
  wire [9:0] _T_29296;
  wire [9:0] _T_29297;
  wire  _T_29299;
  wire [9:0] _T_29305;
  wire [9:0] _T_29306;
  wire  _T_29308;
  wire [9:0] _T_29314;
  wire [9:0] _T_29315;
  wire  _T_29317;
  wire [9:0] _T_29323;
  wire [9:0] _T_29324;
  wire  _T_29326;
  wire [9:0] _T_29332;
  wire [9:0] _T_29333;
  wire  _T_29335;
  wire [9:0] _T_29341;
  wire [9:0] _T_29342;
  wire  _T_29344;
  wire [9:0] _T_29350;
  wire [9:0] _T_29351;
  wire  _T_29353;
  wire [9:0] _T_29359;
  wire [9:0] _T_29360;
  wire  _T_29362;
  wire [9:0] _T_29368;
  wire [9:0] _T_29369;
  wire  _T_29371;
  wire [9:0] _T_29377;
  wire [9:0] _T_29378;
  wire  _T_29380;
  wire [9:0] _T_29386;
  wire [9:0] _T_29387;
  wire  _T_29389;
  wire [9:0] _T_29395;
  wire [9:0] _T_29396;
  wire  _T_29398;
  wire [9:0] _T_29404;
  wire [9:0] _T_29405;
  wire  _T_29407;
  wire [9:0] _T_29413;
  wire [9:0] _T_29414;
  wire  _T_29416;
  wire [9:0] _T_29422;
  wire [9:0] _T_29423;
  wire  _T_29425;
  wire [9:0] _T_29431;
  wire [9:0] _T_29432;
  wire  _T_29434;
  wire [9:0] _T_29440;
  wire [9:0] _T_29441;
  wire  _T_29443;
  wire [9:0] _T_29449;
  wire [9:0] _T_29450;
  wire  _T_29452;
  wire [9:0] _T_29458;
  wire [9:0] _T_29459;
  wire  _T_29461;
  wire [9:0] _T_29467;
  wire [9:0] _T_29468;
  wire  _T_29470;
  wire [9:0] _T_29476;
  wire [9:0] _T_29477;
  wire  _T_29479;
  wire [9:0] _T_29485;
  wire [9:0] _T_29486;
  wire  _T_29488;
  wire [9:0] _T_29494;
  wire [9:0] _T_29495;
  wire  _T_29497;
  wire [9:0] _T_29503;
  wire [9:0] _T_29504;
  wire  _T_29506;
  wire [9:0] _T_29512;
  wire [9:0] _T_29513;
  wire  _T_29515;
  wire [9:0] _T_29521;
  wire [9:0] _T_29522;
  wire  _T_29524;
  wire [9:0] _T_29530;
  wire [9:0] _T_29531;
  wire  _T_29533;
  wire [9:0] _T_29539;
  wire [9:0] _T_29540;
  wire  _T_29542;
  wire [9:0] _T_29548;
  wire [9:0] _T_29549;
  wire  _T_29551;
  wire [9:0] _T_29557;
  wire [9:0] _T_29558;
  wire  _T_29560;
  wire [9:0] _T_29566;
  wire [9:0] _T_29567;
  wire  _T_29569;
  wire [9:0] _T_29575;
  wire [9:0] _T_29576;
  wire  _T_29578;
  wire [9:0] _T_29584;
  wire [9:0] _T_29585;
  wire  _T_29587;
  wire [9:0] _T_29593;
  wire [9:0] _T_29594;
  wire  _T_29596;
  wire [9:0] _T_29602;
  wire [9:0] _T_29603;
  wire  _T_29605;
  wire [9:0] _T_29611;
  wire [9:0] _T_29612;
  wire  _T_29614;
  wire [9:0] _T_29620;
  wire [9:0] _T_29621;
  wire  _T_29623;
  wire [9:0] _T_29629;
  wire [9:0] _T_29630;
  wire  _T_29632;
  wire [9:0] _T_29638;
  wire [9:0] _T_29639;
  wire  _T_29641;
  wire [9:0] _T_29647;
  wire [9:0] _T_29648;
  wire  _T_29650;
  wire [9:0] _T_29656;
  wire [9:0] _T_29657;
  wire  _T_29659;
  wire [9:0] _T_29665;
  wire [9:0] _T_29666;
  wire  _T_29668;
  wire [9:0] _T_29674;
  wire [9:0] _T_29675;
  wire  _T_29677;
  wire  _T_34998;
  wire  _T_34999;
  wire  _T_35000;
  wire  _T_35001;
  wire [7:0] _T_35005;
  wire [7:0] _T_35009;
  wire [7:0] _T_35013;
  wire [7:0] _T_35017;
  wire [15:0] _T_35018;
  wire [15:0] _T_35019;
  wire [31:0] _T_35020;
  wire [7:0] _T_35044;
  wire [7:0] _T_35048;
  wire  _T_35050;
  wire [7:0] _T_35064;
  wire [7:0] _T_35084;
  wire [7:0] _T_35088;
  wire  _T_35090;
  wire [7:0] _T_35104;
  wire [15:0] _GEN_5773;
  wire [15:0] _T_35119;
  wire [15:0] _GEN_5774;
  wire [15:0] _T_35123;
  wire [7:0] _T_35124;
  wire [7:0] _T_35128;
  wire  _T_35130;
  wire [7:0] _T_35144;
  wire [23:0] _GEN_5775;
  wire [23:0] _T_35159;
  wire [23:0] _GEN_5776;
  wire [23:0] _T_35163;
  wire [7:0] _T_35164;
  wire [7:0] _T_35168;
  wire  _T_35170;
  wire [7:0] _T_35184;
  wire [31:0] _GEN_5777;
  wire [31:0] _T_35199;
  wire [31:0] _GEN_5778;
  wire [31:0] _T_35203;
  wire [15:0] _GEN_5779;
  wire [15:0] _T_35279;
  wire [15:0] _GEN_5780;
  wire [15:0] _T_35283;
  wire [23:0] _GEN_5781;
  wire [23:0] _T_35319;
  wire [23:0] _GEN_5782;
  wire [23:0] _T_35323;
  wire [31:0] _GEN_5783;
  wire [31:0] _T_35359;
  wire [31:0] _GEN_5784;
  wire [31:0] _T_35363;
  wire [15:0] _GEN_5785;
  wire [15:0] _T_35439;
  wire [15:0] _GEN_5786;
  wire [15:0] _T_35443;
  wire [23:0] _GEN_5787;
  wire [23:0] _T_35479;
  wire [23:0] _GEN_5788;
  wire [23:0] _T_35483;
  wire [31:0] _GEN_5789;
  wire [31:0] _T_35519;
  wire [31:0] _GEN_5790;
  wire [31:0] _T_35523;
  wire [15:0] _GEN_5791;
  wire [15:0] _T_35599;
  wire [15:0] _GEN_5792;
  wire [15:0] _T_35603;
  wire [23:0] _GEN_5793;
  wire [23:0] _T_35639;
  wire [23:0] _GEN_5794;
  wire [23:0] _T_35643;
  wire [31:0] _GEN_5795;
  wire [31:0] _T_35679;
  wire [31:0] _GEN_5796;
  wire [31:0] _T_35683;
  wire [15:0] _GEN_5797;
  wire [15:0] _T_35919;
  wire [15:0] _GEN_5798;
  wire [15:0] _T_35923;
  wire [23:0] _GEN_5799;
  wire [23:0] _T_35959;
  wire [23:0] _GEN_5800;
  wire [23:0] _T_35963;
  wire [31:0] _GEN_5801;
  wire [31:0] _T_35999;
  wire [31:0] _GEN_5802;
  wire [31:0] _T_36003;
  wire [15:0] _GEN_5803;
  wire [15:0] _T_36079;
  wire [15:0] _GEN_5804;
  wire [15:0] _T_36083;
  wire [23:0] _GEN_5805;
  wire [23:0] _T_36119;
  wire [23:0] _GEN_5806;
  wire [23:0] _T_36123;
  wire [31:0] _GEN_5807;
  wire [31:0] _T_36159;
  wire [31:0] _GEN_5808;
  wire [31:0] _T_36163;
  wire [15:0] _GEN_5809;
  wire [15:0] _T_36239;
  wire [15:0] _GEN_5810;
  wire [15:0] _T_36243;
  wire [23:0] _GEN_5811;
  wire [23:0] _T_36279;
  wire [23:0] _GEN_5812;
  wire [23:0] _T_36283;
  wire [31:0] _GEN_5813;
  wire [31:0] _T_36319;
  wire [31:0] _GEN_5814;
  wire [31:0] _T_36323;
  wire [15:0] _GEN_5815;
  wire [15:0] _T_36399;
  wire [15:0] _GEN_5816;
  wire [15:0] _T_36403;
  wire [23:0] _GEN_5817;
  wire [23:0] _T_36439;
  wire [23:0] _GEN_5818;
  wire [23:0] _T_36443;
  wire [31:0] _GEN_5819;
  wire [31:0] _T_36479;
  wire [31:0] _GEN_5820;
  wire [31:0] _T_36483;
  wire  _T_36663;
  wire [7:0] _GEN_2439;
  wire  _T_36703;
  wire [7:0] _GEN_2440;
  wire  _T_36743;
  wire [7:0] _GEN_2441;
  wire  _T_36783;
  wire [7:0] _GEN_2442;
  wire [15:0] _GEN_5827;
  wire [15:0] _T_36879;
  wire [15:0] _GEN_5828;
  wire [15:0] _T_36883;
  wire [23:0] _GEN_5829;
  wire [23:0] _T_36919;
  wire [23:0] _GEN_5830;
  wire [23:0] _T_36923;
  wire [31:0] _GEN_5831;
  wire [31:0] _T_36959;
  wire [31:0] _GEN_5832;
  wire [31:0] _T_36963;
  wire [15:0] _GEN_5833;
  wire [15:0] _T_37039;
  wire [15:0] _GEN_5834;
  wire [15:0] _T_37043;
  wire [23:0] _GEN_5835;
  wire [23:0] _T_37079;
  wire [23:0] _GEN_5836;
  wire [23:0] _T_37083;
  wire [31:0] _GEN_5837;
  wire [31:0] _T_37119;
  wire [31:0] _GEN_5838;
  wire [31:0] _T_37123;
  wire [15:0] _GEN_5839;
  wire [15:0] _T_37199;
  wire [15:0] _GEN_5840;
  wire [15:0] _T_37203;
  wire [23:0] _GEN_5841;
  wire [23:0] _T_37239;
  wire [23:0] _GEN_5842;
  wire [23:0] _T_37243;
  wire [31:0] _GEN_5843;
  wire [31:0] _T_37279;
  wire [31:0] _GEN_5844;
  wire [31:0] _T_37283;
  wire [15:0] _GEN_5845;
  wire [15:0] _T_37359;
  wire [15:0] _GEN_5846;
  wire [15:0] _T_37363;
  wire [23:0] _GEN_5847;
  wire [23:0] _T_37399;
  wire [23:0] _GEN_5848;
  wire [23:0] _T_37403;
  wire [31:0] _GEN_5849;
  wire [31:0] _T_37439;
  wire [31:0] _GEN_5850;
  wire [31:0] _T_37443;
  wire [15:0] _GEN_5851;
  wire [15:0] _T_37519;
  wire [15:0] _GEN_5852;
  wire [15:0] _T_37523;
  wire [23:0] _GEN_5853;
  wire [23:0] _T_37559;
  wire [23:0] _GEN_5854;
  wire [23:0] _T_37563;
  wire [31:0] _GEN_5855;
  wire [31:0] _T_37599;
  wire [31:0] _GEN_5856;
  wire [31:0] _T_37603;
  wire [15:0] _GEN_5857;
  wire [15:0] _T_37679;
  wire [15:0] _GEN_5858;
  wire [15:0] _T_37683;
  wire [23:0] _GEN_5859;
  wire [23:0] _T_37719;
  wire [23:0] _GEN_5860;
  wire [23:0] _T_37723;
  wire [31:0] _GEN_5861;
  wire [31:0] _T_37759;
  wire [31:0] _GEN_5862;
  wire [31:0] _T_37763;
  wire [15:0] _GEN_5863;
  wire [15:0] _T_37839;
  wire [15:0] _GEN_5864;
  wire [15:0] _T_37843;
  wire [23:0] _GEN_5865;
  wire [23:0] _T_37879;
  wire [23:0] _GEN_5866;
  wire [23:0] _T_37883;
  wire [31:0] _GEN_5867;
  wire [31:0] _T_37919;
  wire [31:0] _GEN_5868;
  wire [31:0] _T_37923;
  wire [15:0] _GEN_5869;
  wire [15:0] _T_37999;
  wire [15:0] _GEN_5870;
  wire [15:0] _T_38003;
  wire [23:0] _GEN_5871;
  wire [23:0] _T_38039;
  wire [23:0] _GEN_5872;
  wire [23:0] _T_38043;
  wire [31:0] _GEN_5873;
  wire [31:0] _T_38079;
  wire [31:0] _GEN_5874;
  wire [31:0] _T_38083;
  wire [15:0] _GEN_5875;
  wire [15:0] _T_38159;
  wire [15:0] _GEN_5876;
  wire [15:0] _T_38163;
  wire [23:0] _GEN_5877;
  wire [23:0] _T_38199;
  wire [23:0] _GEN_5878;
  wire [23:0] _T_38203;
  wire [31:0] _GEN_5879;
  wire [31:0] _T_38239;
  wire [31:0] _GEN_5880;
  wire [31:0] _T_38243;
  wire [15:0] _GEN_5881;
  wire [15:0] _T_38479;
  wire [15:0] _GEN_5882;
  wire [15:0] _T_38483;
  wire [23:0] _GEN_5883;
  wire [23:0] _T_38519;
  wire [23:0] _GEN_5884;
  wire [23:0] _T_38523;
  wire [31:0] _GEN_5885;
  wire [31:0] _T_38559;
  wire [31:0] _GEN_5886;
  wire [31:0] _T_38563;
  wire [15:0] _GEN_5887;
  wire [15:0] _T_38639;
  wire [15:0] _GEN_5888;
  wire [15:0] _T_38643;
  wire [23:0] _GEN_5889;
  wire [23:0] _T_38679;
  wire [23:0] _GEN_5890;
  wire [23:0] _T_38683;
  wire [31:0] _GEN_5891;
  wire [31:0] _T_38719;
  wire [31:0] _GEN_5892;
  wire [31:0] _T_38723;
  wire [15:0] _GEN_5893;
  wire [15:0] _T_38799;
  wire [15:0] _GEN_5894;
  wire [15:0] _T_38803;
  wire [23:0] _GEN_5895;
  wire [23:0] _T_38839;
  wire [23:0] _GEN_5896;
  wire [23:0] _T_38843;
  wire [31:0] _GEN_5897;
  wire [31:0] _T_38879;
  wire [31:0] _GEN_5898;
  wire [31:0] _T_38883;
  wire [15:0] _GEN_5899;
  wire [15:0] _T_38959;
  wire [15:0] _GEN_5900;
  wire [15:0] _T_38963;
  wire [23:0] _GEN_5901;
  wire [23:0] _T_38999;
  wire [23:0] _GEN_5902;
  wire [23:0] _T_39003;
  wire [31:0] _GEN_5903;
  wire [31:0] _T_39039;
  wire [31:0] _GEN_5904;
  wire [31:0] _T_39043;
  wire [15:0] _GEN_5905;
  wire [15:0] _T_39119;
  wire [15:0] _GEN_5906;
  wire [15:0] _T_39123;
  wire [23:0] _GEN_5907;
  wire [23:0] _T_39159;
  wire [23:0] _GEN_5908;
  wire [23:0] _T_39163;
  wire [31:0] _GEN_5909;
  wire [31:0] _T_39199;
  wire [31:0] _GEN_5910;
  wire [31:0] _T_39203;
  wire [15:0] _GEN_5911;
  wire [15:0] _T_39279;
  wire [15:0] _GEN_5912;
  wire [15:0] _T_39283;
  wire [23:0] _GEN_5913;
  wire [23:0] _T_39319;
  wire [23:0] _GEN_5914;
  wire [23:0] _T_39323;
  wire [31:0] _GEN_5915;
  wire [31:0] _T_39359;
  wire [31:0] _GEN_5916;
  wire [31:0] _T_39363;
  wire [15:0] _GEN_5917;
  wire [15:0] _T_39439;
  wire [15:0] _GEN_5918;
  wire [15:0] _T_39443;
  wire [23:0] _GEN_5919;
  wire [23:0] _T_39479;
  wire [23:0] _GEN_5920;
  wire [23:0] _T_39483;
  wire [31:0] _GEN_5921;
  wire [31:0] _T_39519;
  wire [31:0] _GEN_5922;
  wire [31:0] _T_39523;
  wire [15:0] _GEN_5923;
  wire [15:0] _T_39599;
  wire [15:0] _GEN_5924;
  wire [15:0] _T_39603;
  wire [23:0] _GEN_5925;
  wire [23:0] _T_39639;
  wire [23:0] _GEN_5926;
  wire [23:0] _T_39643;
  wire [31:0] _GEN_5927;
  wire [31:0] _T_39679;
  wire [31:0] _GEN_5928;
  wire [31:0] _T_39683;
  wire [15:0] _GEN_5929;
  wire [15:0] _T_39759;
  wire [15:0] _GEN_5930;
  wire [15:0] _T_39763;
  wire [23:0] _GEN_5931;
  wire [23:0] _T_39799;
  wire [23:0] _GEN_5932;
  wire [23:0] _T_39803;
  wire [31:0] _GEN_5933;
  wire [31:0] _T_39839;
  wire [31:0] _GEN_5934;
  wire [31:0] _T_39843;
  wire [15:0] _GEN_5935;
  wire [15:0] _T_39919;
  wire [15:0] _GEN_5936;
  wire [15:0] _T_39923;
  wire [23:0] _GEN_5937;
  wire [23:0] _T_39959;
  wire [23:0] _GEN_5938;
  wire [23:0] _T_39963;
  wire [31:0] _GEN_5939;
  wire [31:0] _T_39999;
  wire [31:0] _GEN_5940;
  wire [31:0] _T_40003;
  wire [15:0] _GEN_5941;
  wire [15:0] _T_40079;
  wire [15:0] _GEN_5942;
  wire [15:0] _T_40083;
  wire [23:0] _GEN_5943;
  wire [23:0] _T_40119;
  wire [23:0] _GEN_5944;
  wire [23:0] _T_40123;
  wire [31:0] _GEN_5945;
  wire [31:0] _T_40159;
  wire [31:0] _GEN_5946;
  wire [31:0] _T_40163;
  wire [15:0] _GEN_5947;
  wire [15:0] _T_40239;
  wire [15:0] _GEN_5948;
  wire [15:0] _T_40243;
  wire [23:0] _GEN_5949;
  wire [23:0] _T_40279;
  wire [23:0] _GEN_5950;
  wire [23:0] _T_40283;
  wire [31:0] _GEN_5951;
  wire [31:0] _T_40319;
  wire [31:0] _GEN_5952;
  wire [31:0] _T_40323;
  wire [15:0] _GEN_5953;
  wire [15:0] _T_40399;
  wire [15:0] _GEN_5954;
  wire [15:0] _T_40403;
  wire [23:0] _GEN_5955;
  wire [23:0] _T_40439;
  wire [23:0] _GEN_5956;
  wire [23:0] _T_40443;
  wire [31:0] _GEN_5957;
  wire [31:0] _T_40479;
  wire [31:0] _GEN_5958;
  wire [31:0] _T_40483;
  wire [15:0] _GEN_5959;
  wire [15:0] _T_40559;
  wire [15:0] _GEN_5960;
  wire [15:0] _T_40563;
  wire [23:0] _GEN_5961;
  wire [23:0] _T_40599;
  wire [23:0] _GEN_5962;
  wire [23:0] _T_40603;
  wire [31:0] _GEN_5963;
  wire [31:0] _T_40639;
  wire [31:0] _GEN_5964;
  wire [31:0] _T_40643;
  wire [15:0] _GEN_5965;
  wire [15:0] _T_40719;
  wire [15:0] _GEN_5966;
  wire [15:0] _T_40723;
  wire [23:0] _GEN_5967;
  wire [23:0] _T_40759;
  wire [23:0] _GEN_5968;
  wire [23:0] _T_40763;
  wire [31:0] _GEN_5969;
  wire [31:0] _T_40799;
  wire [31:0] _GEN_5970;
  wire [31:0] _T_40803;
  wire [15:0] _GEN_5971;
  wire [15:0] _T_40879;
  wire [15:0] _GEN_5972;
  wire [15:0] _T_40883;
  wire [23:0] _GEN_5973;
  wire [23:0] _T_40919;
  wire [23:0] _GEN_5974;
  wire [23:0] _T_40923;
  wire [31:0] _GEN_5975;
  wire [31:0] _T_40959;
  wire [31:0] _GEN_5976;
  wire [31:0] _T_40963;
  wire [15:0] _GEN_5977;
  wire [15:0] _T_41039;
  wire [15:0] _GEN_5978;
  wire [15:0] _T_41043;
  wire [23:0] _GEN_5979;
  wire [23:0] _T_41079;
  wire [23:0] _GEN_5980;
  wire [23:0] _T_41083;
  wire [31:0] _GEN_5981;
  wire [31:0] _T_41119;
  wire [31:0] _GEN_5982;
  wire [31:0] _T_41123;
  wire [15:0] _GEN_5983;
  wire [15:0] _T_41199;
  wire [15:0] _GEN_5984;
  wire [15:0] _T_41203;
  wire [23:0] _GEN_5985;
  wire [23:0] _T_41239;
  wire [23:0] _GEN_5986;
  wire [23:0] _T_41243;
  wire [31:0] _GEN_5987;
  wire [31:0] _T_41279;
  wire [31:0] _GEN_5988;
  wire [31:0] _T_41283;
  wire [15:0] _GEN_5989;
  wire [15:0] _T_41359;
  wire [15:0] _GEN_5990;
  wire [15:0] _T_41363;
  wire [23:0] _GEN_5991;
  wire [23:0] _T_41399;
  wire [23:0] _GEN_5992;
  wire [23:0] _T_41403;
  wire [31:0] _GEN_5993;
  wire [31:0] _T_41439;
  wire [31:0] _GEN_5994;
  wire [31:0] _T_41443;
  wire [15:0] _GEN_5995;
  wire [15:0] _T_41519;
  wire [15:0] _GEN_5996;
  wire [15:0] _T_41523;
  wire [23:0] _GEN_5997;
  wire [23:0] _T_41559;
  wire [23:0] _GEN_5998;
  wire [23:0] _T_41563;
  wire [31:0] _GEN_5999;
  wire [31:0] _T_41599;
  wire [31:0] _GEN_6000;
  wire [31:0] _T_41603;
  wire [15:0] _GEN_6001;
  wire [15:0] _T_41679;
  wire [15:0] _GEN_6002;
  wire [15:0] _T_41683;
  wire [23:0] _GEN_6003;
  wire [23:0] _T_41719;
  wire [23:0] _GEN_6004;
  wire [23:0] _T_41723;
  wire [31:0] _GEN_6005;
  wire [31:0] _T_41759;
  wire [31:0] _GEN_6006;
  wire [31:0] _T_41763;
  wire [15:0] _GEN_6007;
  wire [15:0] _T_41839;
  wire [15:0] _GEN_6008;
  wire [15:0] _T_41843;
  wire [23:0] _GEN_6009;
  wire [23:0] _T_41879;
  wire [23:0] _GEN_6010;
  wire [23:0] _T_41883;
  wire [31:0] _GEN_6011;
  wire [31:0] _T_41919;
  wire [31:0] _GEN_6012;
  wire [31:0] _T_41923;
  wire [15:0] _GEN_6013;
  wire [15:0] _T_41999;
  wire [15:0] _GEN_6014;
  wire [15:0] _T_42003;
  wire [23:0] _GEN_6015;
  wire [23:0] _T_42039;
  wire [23:0] _GEN_6016;
  wire [23:0] _T_42043;
  wire [31:0] _GEN_6017;
  wire [31:0] _T_42079;
  wire [31:0] _GEN_6018;
  wire [31:0] _T_42083;
  wire [15:0] _GEN_6019;
  wire [15:0] _T_42159;
  wire [15:0] _GEN_6020;
  wire [15:0] _T_42163;
  wire [23:0] _GEN_6021;
  wire [23:0] _T_42199;
  wire [23:0] _GEN_6022;
  wire [23:0] _T_42203;
  wire [31:0] _GEN_6023;
  wire [31:0] _T_42239;
  wire [31:0] _GEN_6024;
  wire [31:0] _T_42243;
  wire  _T_42263;
  wire [7:0] _GEN_2443;
  wire  _T_42303;
  wire [7:0] _GEN_2444;
  wire  _T_42343;
  wire [7:0] _GEN_2445;
  wire  _T_42383;
  wire [7:0] _GEN_2446;
  wire [15:0] _GEN_6031;
  wire [15:0] _T_42479;
  wire [15:0] _GEN_6032;
  wire [15:0] _T_42483;
  wire [23:0] _GEN_6033;
  wire [23:0] _T_42519;
  wire [23:0] _GEN_6034;
  wire [23:0] _T_42523;
  wire [31:0] _GEN_6035;
  wire [31:0] _T_42559;
  wire [31:0] _GEN_6036;
  wire [31:0] _T_42563;
  wire [15:0] _GEN_6037;
  wire [15:0] _T_42639;
  wire [15:0] _GEN_6038;
  wire [15:0] _T_42643;
  wire [23:0] _GEN_6039;
  wire [23:0] _T_42679;
  wire [23:0] _GEN_6040;
  wire [23:0] _T_42683;
  wire [31:0] _GEN_6041;
  wire [31:0] _T_42719;
  wire [31:0] _GEN_6042;
  wire [31:0] _T_42723;
  wire [15:0] _GEN_6043;
  wire [15:0] _T_42799;
  wire [15:0] _GEN_6044;
  wire [15:0] _T_42803;
  wire [23:0] _GEN_6045;
  wire [23:0] _T_42839;
  wire [23:0] _GEN_6046;
  wire [23:0] _T_42843;
  wire [31:0] _GEN_6047;
  wire [31:0] _T_42879;
  wire [31:0] _GEN_6048;
  wire [31:0] _T_42883;
  wire [15:0] _GEN_6049;
  wire [15:0] _T_42959;
  wire [15:0] _GEN_6050;
  wire [15:0] _T_42963;
  wire [23:0] _GEN_6051;
  wire [23:0] _T_42999;
  wire [23:0] _GEN_6052;
  wire [23:0] _T_43003;
  wire [31:0] _GEN_6053;
  wire [31:0] _T_43039;
  wire [31:0] _GEN_6054;
  wire [31:0] _T_43043;
  wire [15:0] _GEN_6055;
  wire [15:0] _T_43119;
  wire [15:0] _GEN_6056;
  wire [15:0] _T_43123;
  wire [23:0] _GEN_6057;
  wire [23:0] _T_43159;
  wire [23:0] _GEN_6058;
  wire [23:0] _T_43163;
  wire [31:0] _GEN_6059;
  wire [31:0] _T_43199;
  wire [31:0] _GEN_6060;
  wire [31:0] _T_43203;
  wire  _T_43223;
  wire [7:0] _GEN_2447;
  wire  _T_43263;
  wire [7:0] _GEN_2448;
  wire  _T_43303;
  wire [7:0] _GEN_2449;
  wire  _T_43343;
  wire [7:0] _GEN_2450;
  wire [15:0] _GEN_6067;
  wire [15:0] _T_43439;
  wire [15:0] _GEN_6068;
  wire [15:0] _T_43443;
  wire [23:0] _GEN_6069;
  wire [23:0] _T_43479;
  wire [23:0] _GEN_6070;
  wire [23:0] _T_43483;
  wire [31:0] _GEN_6071;
  wire [31:0] _T_43519;
  wire [31:0] _GEN_6072;
  wire [31:0] _T_43523;
  wire [15:0] _GEN_6073;
  wire [15:0] _T_43759;
  wire [15:0] _GEN_6074;
  wire [15:0] _T_43763;
  wire [23:0] _GEN_6075;
  wire [23:0] _T_43799;
  wire [23:0] _GEN_6076;
  wire [23:0] _T_43803;
  wire [31:0] _GEN_6077;
  wire [31:0] _T_43839;
  wire [31:0] _GEN_6078;
  wire [31:0] _T_43843;
  wire [15:0] _GEN_6079;
  wire [15:0] _T_43919;
  wire [15:0] _GEN_6080;
  wire [15:0] _T_43923;
  wire [23:0] _GEN_6081;
  wire [23:0] _T_43959;
  wire [23:0] _GEN_6082;
  wire [23:0] _T_43963;
  wire [31:0] _GEN_6083;
  wire [31:0] _T_43999;
  wire [31:0] _GEN_6084;
  wire [31:0] _T_44003;
  wire [15:0] _GEN_6085;
  wire [15:0] _T_44079;
  wire [15:0] _GEN_6086;
  wire [15:0] _T_44083;
  wire [23:0] _GEN_6087;
  wire [23:0] _T_44119;
  wire [23:0] _GEN_6088;
  wire [23:0] _T_44123;
  wire [31:0] _GEN_6089;
  wire [31:0] _T_44159;
  wire [31:0] _GEN_6090;
  wire [31:0] _T_44163;
  wire [15:0] _GEN_6091;
  wire [15:0] _T_44239;
  wire [15:0] _GEN_6092;
  wire [15:0] _T_44243;
  wire [23:0] _GEN_6093;
  wire [23:0] _T_44279;
  wire [23:0] _GEN_6094;
  wire [23:0] _T_44283;
  wire [31:0] _GEN_6095;
  wire [31:0] _T_44319;
  wire [31:0] _GEN_6096;
  wire [31:0] _T_44323;
  wire [15:0] _GEN_6097;
  wire [15:0] _T_44399;
  wire [15:0] _GEN_6098;
  wire [15:0] _T_44403;
  wire [23:0] _GEN_6099;
  wire [23:0] _T_44439;
  wire [23:0] _GEN_6100;
  wire [23:0] _T_44443;
  wire [31:0] _GEN_6101;
  wire [31:0] _T_44479;
  wire [31:0] _GEN_6102;
  wire [31:0] _T_44483;
  wire  _T_44503;
  wire [7:0] _GEN_2451;
  wire  _T_44543;
  wire [7:0] _GEN_2452;
  wire  _T_44583;
  wire [7:0] _GEN_2453;
  wire  _T_44623;
  wire [7:0] _GEN_2454;
  wire [15:0] _GEN_6109;
  wire [15:0] _T_44719;
  wire [15:0] _GEN_6110;
  wire [15:0] _T_44723;
  wire [23:0] _GEN_6111;
  wire [23:0] _T_44759;
  wire [23:0] _GEN_6112;
  wire [23:0] _T_44763;
  wire [31:0] _GEN_6113;
  wire [31:0] _T_44799;
  wire [31:0] _GEN_6114;
  wire [31:0] _T_44803;
  wire [15:0] _GEN_6115;
  wire [15:0] _T_44879;
  wire [15:0] _GEN_6116;
  wire [15:0] _T_44883;
  wire [23:0] _GEN_6117;
  wire [23:0] _T_44919;
  wire [23:0] _GEN_6118;
  wire [23:0] _T_44923;
  wire [31:0] _GEN_6119;
  wire [31:0] _T_44959;
  wire [31:0] _GEN_6120;
  wire [31:0] _T_44963;
  wire [15:0] _GEN_6121;
  wire [15:0] _T_45039;
  wire [15:0] _GEN_6122;
  wire [15:0] _T_45043;
  wire [23:0] _GEN_6123;
  wire [23:0] _T_45079;
  wire [23:0] _GEN_6124;
  wire [23:0] _T_45083;
  wire [31:0] _GEN_6125;
  wire [31:0] _T_45119;
  wire [31:0] _GEN_6126;
  wire [31:0] _T_45123;
  wire [15:0] _GEN_6127;
  wire [15:0] _T_45199;
  wire [15:0] _GEN_6128;
  wire [15:0] _T_45203;
  wire [23:0] _GEN_6129;
  wire [23:0] _T_45239;
  wire [23:0] _GEN_6130;
  wire [23:0] _T_45243;
  wire [31:0] _GEN_6131;
  wire [31:0] _T_45279;
  wire [31:0] _GEN_6132;
  wire [31:0] _T_45283;
  wire [15:0] _GEN_6133;
  wire [15:0] _T_45359;
  wire [15:0] _GEN_6134;
  wire [15:0] _T_45363;
  wire [23:0] _GEN_6135;
  wire [23:0] _T_45399;
  wire [23:0] _GEN_6136;
  wire [23:0] _T_45403;
  wire [31:0] _GEN_6137;
  wire [31:0] _T_45439;
  wire [31:0] _GEN_6138;
  wire [31:0] _T_45443;
  wire [15:0] _GEN_6139;
  wire [15:0] _T_45519;
  wire [15:0] _GEN_6140;
  wire [15:0] _T_45523;
  wire [23:0] _GEN_6141;
  wire [23:0] _T_45559;
  wire [23:0] _GEN_6142;
  wire [23:0] _T_45563;
  wire [31:0] _GEN_6143;
  wire [31:0] _T_45599;
  wire [31:0] _GEN_6144;
  wire [31:0] _T_45603;
  wire [15:0] _GEN_6145;
  wire [15:0] _T_45679;
  wire [15:0] _GEN_6146;
  wire [15:0] _T_45683;
  wire [23:0] _GEN_6147;
  wire [23:0] _T_45719;
  wire [23:0] _GEN_6148;
  wire [23:0] _T_45723;
  wire [31:0] _GEN_6149;
  wire [31:0] _T_45759;
  wire [31:0] _GEN_6150;
  wire [31:0] _T_45763;
  wire [15:0] _GEN_6151;
  wire [15:0] _T_45999;
  wire [15:0] _GEN_6152;
  wire [15:0] _T_46003;
  wire [23:0] _GEN_6153;
  wire [23:0] _T_46039;
  wire [23:0] _GEN_6154;
  wire [23:0] _T_46043;
  wire [31:0] _GEN_6155;
  wire [31:0] _T_46079;
  wire [31:0] _GEN_6156;
  wire [31:0] _T_46083;
  wire [15:0] _GEN_6157;
  wire [15:0] _T_46199;
  wire [15:0] _GEN_6158;
  wire [15:0] _T_46203;
  wire [23:0] _GEN_6159;
  wire [23:0] _T_46239;
  wire [23:0] _GEN_6160;
  wire [23:0] _T_46243;
  wire [31:0] _GEN_6161;
  wire [31:0] _T_46279;
  wire [31:0] _GEN_6162;
  wire [31:0] _T_46283;
  wire [15:0] _GEN_6163;
  wire [15:0] _T_46359;
  wire [15:0] _GEN_6164;
  wire [15:0] _T_46363;
  wire [23:0] _GEN_6165;
  wire [23:0] _T_46399;
  wire [23:0] _GEN_6166;
  wire [23:0] _T_46403;
  wire [31:0] _GEN_6167;
  wire [31:0] _T_46439;
  wire [31:0] _GEN_6168;
  wire [31:0] _T_46443;
  wire [15:0] _GEN_6169;
  wire [15:0] _T_46519;
  wire [15:0] _GEN_6170;
  wire [15:0] _T_46523;
  wire [23:0] _GEN_6171;
  wire [23:0] _T_46559;
  wire [23:0] _GEN_6172;
  wire [23:0] _T_46563;
  wire [31:0] _GEN_6173;
  wire [31:0] _T_46599;
  wire [31:0] _GEN_6174;
  wire [31:0] _T_46603;
  wire [15:0] _GEN_6175;
  wire [15:0] _T_46679;
  wire [15:0] _GEN_6176;
  wire [15:0] _T_46683;
  wire [23:0] _GEN_6177;
  wire [23:0] _T_46719;
  wire [23:0] _GEN_6178;
  wire [23:0] _T_46723;
  wire [31:0] _GEN_6179;
  wire [31:0] _T_46759;
  wire [31:0] _GEN_6180;
  wire [31:0] _T_46763;
  wire [15:0] _GEN_6181;
  wire [15:0] _T_46999;
  wire [15:0] _GEN_6182;
  wire [15:0] _T_47003;
  wire [23:0] _GEN_6183;
  wire [23:0] _T_47039;
  wire [23:0] _GEN_6184;
  wire [23:0] _T_47043;
  wire [31:0] _GEN_6185;
  wire [31:0] _T_47079;
  wire [31:0] _GEN_6186;
  wire [31:0] _T_47083;
  wire [15:0] _GEN_6187;
  wire [15:0] _T_47159;
  wire [15:0] _GEN_6188;
  wire [15:0] _T_47163;
  wire [23:0] _GEN_6189;
  wire [23:0] _T_47199;
  wire [23:0] _GEN_6190;
  wire [23:0] _T_47203;
  wire [31:0] _GEN_6191;
  wire [31:0] _T_47239;
  wire [31:0] _GEN_6192;
  wire [31:0] _T_47243;
  wire [15:0] _GEN_6193;
  wire [15:0] _T_47479;
  wire [15:0] _GEN_6194;
  wire [15:0] _T_47483;
  wire [23:0] _GEN_6195;
  wire [23:0] _T_47519;
  wire [23:0] _GEN_6196;
  wire [23:0] _T_47523;
  wire [31:0] _GEN_6197;
  wire [31:0] _T_47559;
  wire [31:0] _GEN_6198;
  wire [31:0] _T_47563;
  wire  _T_47583;
  wire [7:0] _GEN_2455;
  wire  _T_47623;
  wire [7:0] _GEN_2456;
  wire  _T_47663;
  wire [7:0] _GEN_2457;
  wire  _T_47703;
  wire [7:0] _GEN_2458;
  wire [15:0] _GEN_6205;
  wire [15:0] _T_47799;
  wire [15:0] _GEN_6206;
  wire [15:0] _T_47803;
  wire [23:0] _GEN_6207;
  wire [23:0] _T_47839;
  wire [23:0] _GEN_6208;
  wire [23:0] _T_47843;
  wire [31:0] _GEN_6209;
  wire [31:0] _T_47879;
  wire [31:0] _GEN_6210;
  wire [31:0] _T_47883;
  wire [15:0] _GEN_6211;
  wire [15:0] _T_48119;
  wire [15:0] _GEN_6212;
  wire [15:0] _T_48123;
  wire [23:0] _GEN_6213;
  wire [23:0] _T_48159;
  wire [23:0] _GEN_6214;
  wire [23:0] _T_48163;
  wire [31:0] _GEN_6215;
  wire [31:0] _T_48199;
  wire [31:0] _GEN_6216;
  wire [31:0] _T_48203;
  wire [15:0] _GEN_6217;
  wire [15:0] _T_48279;
  wire [15:0] _GEN_6218;
  wire [15:0] _T_48283;
  wire [23:0] _GEN_6219;
  wire [23:0] _T_48319;
  wire [23:0] _GEN_6220;
  wire [23:0] _T_48323;
  wire [31:0] _GEN_6221;
  wire [31:0] _T_48359;
  wire [31:0] _GEN_6222;
  wire [31:0] _T_48363;
  wire [15:0] _GEN_6223;
  wire [15:0] _T_48439;
  wire [15:0] _GEN_6224;
  wire [15:0] _T_48443;
  wire [23:0] _GEN_6225;
  wire [23:0] _T_48479;
  wire [23:0] _GEN_6226;
  wire [23:0] _T_48483;
  wire [31:0] _GEN_6227;
  wire [31:0] _T_48519;
  wire [31:0] _GEN_6228;
  wire [31:0] _T_48523;
  wire [15:0] _GEN_6229;
  wire [15:0] _T_48599;
  wire [15:0] _GEN_6230;
  wire [15:0] _T_48603;
  wire [23:0] _GEN_6231;
  wire [23:0] _T_48639;
  wire [23:0] _GEN_6232;
  wire [23:0] _T_48643;
  wire [31:0] _GEN_6233;
  wire [31:0] _T_48679;
  wire [31:0] _GEN_6234;
  wire [31:0] _T_48683;
  wire [15:0] _GEN_6235;
  wire [15:0] _T_48759;
  wire [15:0] _GEN_6236;
  wire [15:0] _T_48763;
  wire [23:0] _GEN_6237;
  wire [23:0] _T_48799;
  wire [23:0] _GEN_6238;
  wire [23:0] _T_48803;
  wire [31:0] _GEN_6239;
  wire [31:0] _T_48839;
  wire [31:0] _GEN_6240;
  wire [31:0] _T_48843;
  wire [15:0] _GEN_6241;
  wire [15:0] _T_48919;
  wire [15:0] _GEN_6242;
  wire [15:0] _T_48923;
  wire [23:0] _GEN_6243;
  wire [23:0] _T_48959;
  wire [23:0] _GEN_6244;
  wire [23:0] _T_48963;
  wire [31:0] _GEN_6245;
  wire [31:0] _T_48999;
  wire [31:0] _GEN_6246;
  wire [31:0] _T_49003;
  wire [15:0] _GEN_6247;
  wire [15:0] _T_49079;
  wire [15:0] _GEN_6248;
  wire [15:0] _T_49083;
  wire [23:0] _GEN_6249;
  wire [23:0] _T_49119;
  wire [23:0] _GEN_6250;
  wire [23:0] _T_49123;
  wire [31:0] _GEN_6251;
  wire [31:0] _T_49159;
  wire [31:0] _GEN_6252;
  wire [31:0] _T_49163;
  wire [15:0] _GEN_6253;
  wire [15:0] _T_49279;
  wire [15:0] _GEN_6254;
  wire [15:0] _T_49283;
  wire [23:0] _GEN_6255;
  wire [23:0] _T_49319;
  wire [23:0] _GEN_6256;
  wire [23:0] _T_49323;
  wire [31:0] _GEN_6257;
  wire [31:0] _T_49359;
  wire [31:0] _GEN_6258;
  wire [31:0] _T_49363;
  wire [15:0] _GEN_6259;
  wire [15:0] _T_49439;
  wire [15:0] _GEN_6260;
  wire [15:0] _T_49443;
  wire [23:0] _GEN_6261;
  wire [23:0] _T_49479;
  wire [23:0] _GEN_6262;
  wire [23:0] _T_49483;
  wire [31:0] _GEN_6263;
  wire [31:0] _T_49519;
  wire [31:0] _GEN_6264;
  wire [31:0] _T_49523;
  wire [15:0] _GEN_6265;
  wire [15:0] _T_49599;
  wire [15:0] _GEN_6266;
  wire [15:0] _T_49603;
  wire [23:0] _GEN_6267;
  wire [23:0] _T_49639;
  wire [23:0] _GEN_6268;
  wire [23:0] _T_49643;
  wire [31:0] _GEN_6269;
  wire [31:0] _T_49679;
  wire [31:0] _GEN_6270;
  wire [31:0] _T_49683;
  wire [15:0] _GEN_6271;
  wire [15:0] _T_49759;
  wire [15:0] _GEN_6272;
  wire [15:0] _T_49763;
  wire [23:0] _GEN_6273;
  wire [23:0] _T_49799;
  wire [23:0] _GEN_6274;
  wire [23:0] _T_49803;
  wire [31:0] _GEN_6275;
  wire [31:0] _T_49839;
  wire [31:0] _GEN_6276;
  wire [31:0] _T_49843;
  wire [15:0] _GEN_6277;
  wire [15:0] _T_49919;
  wire [15:0] _GEN_6278;
  wire [15:0] _T_49923;
  wire [23:0] _GEN_6279;
  wire [23:0] _T_49959;
  wire [23:0] _GEN_6280;
  wire [23:0] _T_49963;
  wire [31:0] _GEN_6281;
  wire [31:0] _T_49999;
  wire [31:0] _GEN_6282;
  wire [31:0] _T_50003;
  wire [15:0] _GEN_6283;
  wire [15:0] _T_50079;
  wire [15:0] _GEN_6284;
  wire [15:0] _T_50083;
  wire [23:0] _GEN_6285;
  wire [23:0] _T_50119;
  wire [23:0] _GEN_6286;
  wire [23:0] _T_50123;
  wire [31:0] _GEN_6287;
  wire [31:0] _T_50159;
  wire [31:0] _GEN_6288;
  wire [31:0] _T_50163;
  wire [9:0] _T_50164;
  wire [9:0] _T_50168;
  wire  _T_50170;
  wire  _T_50183;
  wire [9:0] _T_50184;
  wire [15:0] _GEN_6289;
  wire [15:0] _T_50279;
  wire [15:0] _GEN_6290;
  wire [15:0] _T_50283;
  wire [23:0] _GEN_6291;
  wire [23:0] _T_50319;
  wire [23:0] _GEN_6292;
  wire [23:0] _T_50323;
  wire [31:0] _GEN_6293;
  wire [31:0] _T_50359;
  wire [31:0] _GEN_6294;
  wire [31:0] _T_50363;
  wire [15:0] _GEN_6295;
  wire [15:0] _T_50439;
  wire [15:0] _GEN_6296;
  wire [15:0] _T_50443;
  wire [23:0] _GEN_6297;
  wire [23:0] _T_50479;
  wire [23:0] _GEN_6298;
  wire [23:0] _T_50483;
  wire [31:0] _GEN_6299;
  wire [31:0] _T_50519;
  wire [31:0] _GEN_6300;
  wire [31:0] _T_50523;
  wire [15:0] _GEN_6301;
  wire [15:0] _T_50759;
  wire [15:0] _GEN_6302;
  wire [15:0] _T_50763;
  wire [23:0] _GEN_6303;
  wire [23:0] _T_50799;
  wire [23:0] _GEN_6304;
  wire [23:0] _T_50803;
  wire [31:0] _GEN_6305;
  wire [31:0] _T_50839;
  wire [31:0] _GEN_6306;
  wire [31:0] _T_50843;
  wire [15:0] _GEN_6307;
  wire [15:0] _T_50919;
  wire [15:0] _GEN_6308;
  wire [15:0] _T_50923;
  wire [23:0] _GEN_6309;
  wire [23:0] _T_50959;
  wire [23:0] _GEN_6310;
  wire [23:0] _T_50963;
  wire [31:0] _GEN_6311;
  wire [31:0] _T_50999;
  wire [31:0] _GEN_6312;
  wire [31:0] _T_51003;
  wire [15:0] _GEN_6313;
  wire [15:0] _T_51079;
  wire [15:0] _GEN_6314;
  wire [15:0] _T_51083;
  wire [23:0] _GEN_6315;
  wire [23:0] _T_51119;
  wire [23:0] _GEN_6316;
  wire [23:0] _T_51123;
  wire [31:0] _GEN_6317;
  wire [31:0] _T_51159;
  wire [31:0] _GEN_6318;
  wire [31:0] _T_51163;
  wire [15:0] _GEN_6319;
  wire [15:0] _T_51239;
  wire [15:0] _GEN_6320;
  wire [15:0] _T_51243;
  wire [23:0] _GEN_6321;
  wire [23:0] _T_51279;
  wire [23:0] _GEN_6322;
  wire [23:0] _T_51283;
  wire [31:0] _GEN_6323;
  wire [31:0] _T_51319;
  wire [31:0] _GEN_6324;
  wire [31:0] _T_51323;
  wire [15:0] _GEN_6325;
  wire [15:0] _T_51399;
  wire [15:0] _GEN_6326;
  wire [15:0] _T_51403;
  wire [23:0] _GEN_6327;
  wire [23:0] _T_51439;
  wire [23:0] _GEN_6328;
  wire [23:0] _T_51443;
  wire [31:0] _GEN_6329;
  wire [31:0] _T_51479;
  wire [31:0] _GEN_6330;
  wire [31:0] _T_51483;
  wire  _T_51503;
  wire [7:0] _GEN_2460;
  wire  _T_51543;
  wire [7:0] _GEN_2461;
  wire  _T_51583;
  wire [7:0] _GEN_2462;
  wire  _T_51623;
  wire [7:0] _GEN_2463;
  wire [15:0] _GEN_6337;
  wire [15:0] _T_51879;
  wire [15:0] _GEN_6338;
  wire [15:0] _T_51883;
  wire [23:0] _GEN_6339;
  wire [23:0] _T_51919;
  wire [23:0] _GEN_6340;
  wire [23:0] _T_51923;
  wire [31:0] _GEN_6341;
  wire [31:0] _T_51959;
  wire [31:0] _GEN_6342;
  wire [31:0] _T_51963;
  wire [15:0] _GEN_6343;
  wire [15:0] _T_52039;
  wire [15:0] _GEN_6344;
  wire [15:0] _T_52043;
  wire [23:0] _GEN_6345;
  wire [23:0] _T_52079;
  wire [23:0] _GEN_6346;
  wire [23:0] _T_52083;
  wire [31:0] _GEN_6347;
  wire [31:0] _T_52119;
  wire [31:0] _GEN_6348;
  wire [31:0] _T_52123;
  wire [15:0] _GEN_6349;
  wire [15:0] _T_52199;
  wire [15:0] _GEN_6350;
  wire [15:0] _T_52203;
  wire [23:0] _GEN_6351;
  wire [23:0] _T_52239;
  wire [23:0] _GEN_6352;
  wire [23:0] _T_52243;
  wire [31:0] _GEN_6353;
  wire [31:0] _T_52279;
  wire [31:0] _GEN_6354;
  wire [31:0] _T_52283;
  wire [15:0] _GEN_6355;
  wire [15:0] _T_52359;
  wire [15:0] _GEN_6356;
  wire [15:0] _T_52363;
  wire [23:0] _GEN_6357;
  wire [23:0] _T_52399;
  wire [23:0] _GEN_6358;
  wire [23:0] _T_52403;
  wire [31:0] _GEN_6359;
  wire [31:0] _T_52439;
  wire [31:0] _GEN_6360;
  wire [31:0] _T_52443;
  wire [15:0] _GEN_6361;
  wire [15:0] _T_52519;
  wire [15:0] _GEN_6362;
  wire [15:0] _T_52523;
  wire [23:0] _GEN_6363;
  wire [23:0] _T_52559;
  wire [23:0] _GEN_6364;
  wire [23:0] _T_52563;
  wire [31:0] _GEN_6365;
  wire [31:0] _T_52599;
  wire [31:0] _GEN_6366;
  wire [31:0] _T_52603;
  wire [15:0] _GEN_6367;
  wire [15:0] _T_52679;
  wire [15:0] _GEN_6368;
  wire [15:0] _T_52683;
  wire [23:0] _GEN_6369;
  wire [23:0] _T_52719;
  wire [23:0] _GEN_6370;
  wire [23:0] _T_52723;
  wire [31:0] _GEN_6371;
  wire [31:0] _T_52759;
  wire [31:0] _GEN_6372;
  wire [31:0] _T_52763;
  wire [15:0] _GEN_6373;
  wire [15:0] _T_52839;
  wire [15:0] _GEN_6374;
  wire [15:0] _T_52843;
  wire [23:0] _GEN_6375;
  wire [23:0] _T_52879;
  wire [23:0] _GEN_6376;
  wire [23:0] _T_52883;
  wire [31:0] _GEN_6377;
  wire [31:0] _T_52919;
  wire [31:0] _GEN_6378;
  wire [31:0] _T_52923;
  wire [15:0] _GEN_6379;
  wire [15:0] _T_52999;
  wire [15:0] _GEN_6380;
  wire [15:0] _T_53003;
  wire [23:0] _GEN_6381;
  wire [23:0] _T_53039;
  wire [23:0] _GEN_6382;
  wire [23:0] _T_53043;
  wire [31:0] _GEN_6383;
  wire [31:0] _T_53079;
  wire [31:0] _GEN_6384;
  wire [31:0] _T_53083;
  wire [15:0] _GEN_6385;
  wire [15:0] _T_53159;
  wire [15:0] _GEN_6386;
  wire [15:0] _T_53163;
  wire [23:0] _GEN_6387;
  wire [23:0] _T_53199;
  wire [23:0] _GEN_6388;
  wire [23:0] _T_53203;
  wire [31:0] _GEN_6389;
  wire [31:0] _T_53239;
  wire [31:0] _GEN_6390;
  wire [31:0] _T_53243;
  wire [15:0] _GEN_6391;
  wire [15:0] _T_53319;
  wire [15:0] _GEN_6392;
  wire [15:0] _T_53323;
  wire [23:0] _GEN_6393;
  wire [23:0] _T_53359;
  wire [23:0] _GEN_6394;
  wire [23:0] _T_53363;
  wire [31:0] _GEN_6395;
  wire [31:0] _T_53399;
  wire [31:0] _GEN_6396;
  wire [31:0] _T_53403;
  wire [15:0] _GEN_6397;
  wire [15:0] _T_53479;
  wire [15:0] _GEN_6398;
  wire [15:0] _T_53483;
  wire [23:0] _GEN_6399;
  wire [23:0] _T_53519;
  wire [23:0] _GEN_6400;
  wire [23:0] _T_53523;
  wire [31:0] _GEN_6401;
  wire [31:0] _T_53559;
  wire [31:0] _GEN_6402;
  wire [31:0] _T_53563;
  wire [15:0] _GEN_6403;
  wire [15:0] _T_53639;
  wire [15:0] _GEN_6404;
  wire [15:0] _T_53643;
  wire [23:0] _GEN_6405;
  wire [23:0] _T_53679;
  wire [23:0] _GEN_6406;
  wire [23:0] _T_53683;
  wire [31:0] _GEN_6407;
  wire [31:0] _T_53719;
  wire [31:0] _GEN_6408;
  wire [31:0] _T_53723;
  wire [15:0] _GEN_6409;
  wire [15:0] _T_53959;
  wire [15:0] _GEN_6410;
  wire [15:0] _T_53963;
  wire [23:0] _GEN_6411;
  wire [23:0] _T_53999;
  wire [23:0] _GEN_6412;
  wire [23:0] _T_54003;
  wire [31:0] _GEN_6413;
  wire [31:0] _T_54039;
  wire [31:0] _GEN_6414;
  wire [31:0] _T_54043;
  wire  _T_54063;
  wire [7:0] _GEN_2464;
  wire  _T_54103;
  wire [7:0] _GEN_2465;
  wire  _T_54143;
  wire [7:0] _GEN_2466;
  wire  _T_54183;
  wire [7:0] _GEN_2467;
  wire [15:0] _GEN_6421;
  wire [15:0] _T_54279;
  wire [15:0] _GEN_6422;
  wire [15:0] _T_54283;
  wire [23:0] _GEN_6423;
  wire [23:0] _T_54319;
  wire [23:0] _GEN_6424;
  wire [23:0] _T_54323;
  wire [31:0] _GEN_6425;
  wire [31:0] _T_54359;
  wire [31:0] _GEN_6426;
  wire [31:0] _T_54363;
  wire [15:0] _GEN_6427;
  wire [15:0] _T_54599;
  wire [15:0] _GEN_6428;
  wire [15:0] _T_54603;
  wire [23:0] _GEN_6429;
  wire [23:0] _T_54639;
  wire [23:0] _GEN_6430;
  wire [23:0] _T_54643;
  wire [31:0] _GEN_6431;
  wire [31:0] _T_54679;
  wire [31:0] _GEN_6432;
  wire [31:0] _T_54683;
  wire [15:0] _GEN_6433;
  wire [15:0] _T_54759;
  wire [15:0] _GEN_6434;
  wire [15:0] _T_54763;
  wire [23:0] _GEN_6435;
  wire [23:0] _T_54799;
  wire [23:0] _GEN_6436;
  wire [23:0] _T_54803;
  wire [31:0] _GEN_6437;
  wire [31:0] _T_54839;
  wire [31:0] _GEN_6438;
  wire [31:0] _T_54843;
  wire [15:0] _GEN_6439;
  wire [15:0] _T_54919;
  wire [15:0] _GEN_6440;
  wire [15:0] _T_54923;
  wire [23:0] _GEN_6441;
  wire [23:0] _T_54959;
  wire [23:0] _GEN_6442;
  wire [23:0] _T_54963;
  wire [31:0] _GEN_6443;
  wire [31:0] _T_54999;
  wire [31:0] _GEN_6444;
  wire [31:0] _T_55003;
  wire [15:0] _GEN_6445;
  wire [15:0] _T_55079;
  wire [15:0] _GEN_6446;
  wire [15:0] _T_55083;
  wire [23:0] _GEN_6447;
  wire [23:0] _T_55119;
  wire [23:0] _GEN_6448;
  wire [23:0] _T_55123;
  wire [31:0] _GEN_6449;
  wire [31:0] _T_55159;
  wire [31:0] _GEN_6450;
  wire [31:0] _T_55163;
  wire [15:0] _GEN_6451;
  wire [15:0] _T_55239;
  wire [15:0] _GEN_6452;
  wire [15:0] _T_55243;
  wire [23:0] _GEN_6453;
  wire [23:0] _T_55279;
  wire [23:0] _GEN_6454;
  wire [23:0] _T_55283;
  wire [31:0] _GEN_6455;
  wire [31:0] _T_55319;
  wire [31:0] _GEN_6456;
  wire [31:0] _T_55323;
  wire [15:0] _GEN_6457;
  wire [15:0] _T_55399;
  wire [15:0] _GEN_6458;
  wire [15:0] _T_55403;
  wire [23:0] _GEN_6459;
  wire [23:0] _T_55439;
  wire [23:0] _GEN_6460;
  wire [23:0] _T_55443;
  wire [31:0] _GEN_6461;
  wire [31:0] _T_55479;
  wire [31:0] _GEN_6462;
  wire [31:0] _T_55483;
  wire [15:0] _GEN_6463;
  wire [15:0] _T_55559;
  wire [15:0] _GEN_6464;
  wire [15:0] _T_55563;
  wire [23:0] _GEN_6465;
  wire [23:0] _T_55599;
  wire [23:0] _GEN_6466;
  wire [23:0] _T_55603;
  wire [31:0] _GEN_6467;
  wire [31:0] _T_55639;
  wire [31:0] _GEN_6468;
  wire [31:0] _T_55643;
  wire [15:0] _GEN_6469;
  wire [15:0] _T_55719;
  wire [15:0] _GEN_6470;
  wire [15:0] _T_55723;
  wire [23:0] _GEN_6471;
  wire [23:0] _T_55759;
  wire [23:0] _GEN_6472;
  wire [23:0] _T_55763;
  wire [31:0] _GEN_6473;
  wire [31:0] _T_55799;
  wire [31:0] _GEN_6474;
  wire [31:0] _T_55803;
  wire [15:0] _GEN_6475;
  wire [15:0] _T_55879;
  wire [15:0] _GEN_6476;
  wire [15:0] _T_55883;
  wire [23:0] _GEN_6477;
  wire [23:0] _T_55919;
  wire [23:0] _GEN_6478;
  wire [23:0] _T_55923;
  wire [31:0] _GEN_6479;
  wire [31:0] _T_55959;
  wire [31:0] _GEN_6480;
  wire [31:0] _T_55963;
  wire [15:0] _GEN_6481;
  wire [15:0] _T_56199;
  wire [15:0] _GEN_6482;
  wire [15:0] _T_56203;
  wire [23:0] _GEN_6483;
  wire [23:0] _T_56239;
  wire [23:0] _GEN_6484;
  wire [23:0] _T_56243;
  wire [31:0] _GEN_6485;
  wire [31:0] _T_56279;
  wire [31:0] _GEN_6486;
  wire [31:0] _T_56283;
  wire [15:0] _GEN_6487;
  wire [15:0] _T_56359;
  wire [15:0] _GEN_6488;
  wire [15:0] _T_56363;
  wire [23:0] _GEN_6489;
  wire [23:0] _T_56399;
  wire [23:0] _GEN_6490;
  wire [23:0] _T_56403;
  wire [31:0] _GEN_6491;
  wire [31:0] _T_56439;
  wire [31:0] _GEN_6492;
  wire [31:0] _T_56443;
  wire [15:0] _GEN_6493;
  wire [15:0] _T_56519;
  wire [15:0] _GEN_6494;
  wire [15:0] _T_56523;
  wire [23:0] _GEN_6495;
  wire [23:0] _T_56559;
  wire [23:0] _GEN_6496;
  wire [23:0] _T_56563;
  wire [31:0] _GEN_6497;
  wire [31:0] _T_56599;
  wire [31:0] _GEN_6498;
  wire [31:0] _T_56603;
  wire [15:0] _GEN_6499;
  wire [15:0] _T_56839;
  wire [15:0] _GEN_6500;
  wire [15:0] _T_56843;
  wire [23:0] _GEN_6501;
  wire [23:0] _T_56879;
  wire [23:0] _GEN_6502;
  wire [23:0] _T_56883;
  wire [31:0] _GEN_6503;
  wire [31:0] _T_56919;
  wire [31:0] _GEN_6504;
  wire [31:0] _T_56923;
  wire [15:0] _GEN_6505;
  wire [15:0] _T_56999;
  wire [15:0] _GEN_6506;
  wire [15:0] _T_57003;
  wire [23:0] _GEN_6507;
  wire [23:0] _T_57039;
  wire [23:0] _GEN_6508;
  wire [23:0] _T_57043;
  wire [31:0] _GEN_6509;
  wire [31:0] _T_57079;
  wire [31:0] _GEN_6510;
  wire [31:0] _T_57083;
  wire [15:0] _GEN_6511;
  wire [15:0] _T_57159;
  wire [15:0] _GEN_6512;
  wire [15:0] _T_57163;
  wire [23:0] _GEN_6513;
  wire [23:0] _T_57199;
  wire [23:0] _GEN_6514;
  wire [23:0] _T_57203;
  wire [31:0] _GEN_6515;
  wire [31:0] _T_57239;
  wire [31:0] _GEN_6516;
  wire [31:0] _T_57243;
  wire  _T_57263;
  wire [9:0] _T_57264;
  wire [15:0] _GEN_6517;
  wire [15:0] _T_57359;
  wire [15:0] _GEN_6518;
  wire [15:0] _T_57363;
  wire [23:0] _GEN_6519;
  wire [23:0] _T_57399;
  wire [23:0] _GEN_6520;
  wire [23:0] _T_57403;
  wire [31:0] _GEN_6521;
  wire [31:0] _T_57439;
  wire [31:0] _GEN_6522;
  wire [31:0] _T_57443;
  wire [15:0] _GEN_6523;
  wire [15:0] _T_57519;
  wire [15:0] _GEN_6524;
  wire [15:0] _T_57523;
  wire [23:0] _GEN_6525;
  wire [23:0] _T_57559;
  wire [23:0] _GEN_6526;
  wire [23:0] _T_57563;
  wire [31:0] _GEN_6527;
  wire [31:0] _T_57599;
  wire [31:0] _GEN_6528;
  wire [31:0] _T_57603;
  wire [15:0] _GEN_6529;
  wire [15:0] _T_57679;
  wire [15:0] _GEN_6530;
  wire [15:0] _T_57683;
  wire [23:0] _GEN_6531;
  wire [23:0] _T_57719;
  wire [23:0] _GEN_6532;
  wire [23:0] _T_57723;
  wire [31:0] _GEN_6533;
  wire [31:0] _T_57759;
  wire [31:0] _GEN_6534;
  wire [31:0] _T_57763;
  wire [15:0] _GEN_6535;
  wire [15:0] _T_57839;
  wire [15:0] _GEN_6536;
  wire [15:0] _T_57843;
  wire [23:0] _GEN_6537;
  wire [23:0] _T_57879;
  wire [23:0] _GEN_6538;
  wire [23:0] _T_57883;
  wire [31:0] _GEN_6539;
  wire [31:0] _T_57919;
  wire [31:0] _GEN_6540;
  wire [31:0] _T_57923;
  wire [15:0] _GEN_6541;
  wire [15:0] _T_57999;
  wire [15:0] _GEN_6542;
  wire [15:0] _T_58003;
  wire [23:0] _GEN_6543;
  wire [23:0] _T_58039;
  wire [23:0] _GEN_6544;
  wire [23:0] _T_58043;
  wire [31:0] _GEN_6545;
  wire [31:0] _T_58079;
  wire [31:0] _GEN_6546;
  wire [31:0] _T_58083;
  wire [15:0] _GEN_6547;
  wire [15:0] _T_58159;
  wire [15:0] _GEN_6548;
  wire [15:0] _T_58163;
  wire [23:0] _GEN_6549;
  wire [23:0] _T_58199;
  wire [23:0] _GEN_6550;
  wire [23:0] _T_58203;
  wire [31:0] _GEN_6551;
  wire [31:0] _T_58239;
  wire [31:0] _GEN_6552;
  wire [31:0] _T_58243;
  wire [15:0] _GEN_6553;
  wire [15:0] _T_58319;
  wire [15:0] _GEN_6554;
  wire [15:0] _T_58323;
  wire [23:0] _GEN_6555;
  wire [23:0] _T_58359;
  wire [23:0] _GEN_6556;
  wire [23:0] _T_58363;
  wire [31:0] _GEN_6557;
  wire [31:0] _T_58399;
  wire [31:0] _GEN_6558;
  wire [31:0] _T_58403;
  wire [15:0] _GEN_6559;
  wire [15:0] _T_58479;
  wire [15:0] _GEN_6560;
  wire [15:0] _T_58483;
  wire [23:0] _GEN_6561;
  wire [23:0] _T_58519;
  wire [23:0] _GEN_6562;
  wire [23:0] _T_58523;
  wire [31:0] _GEN_6563;
  wire [31:0] _T_58559;
  wire [31:0] _GEN_6564;
  wire [31:0] _T_58563;
  wire [15:0] _GEN_6565;
  wire [15:0] _T_58639;
  wire [15:0] _GEN_6566;
  wire [15:0] _T_58643;
  wire [23:0] _GEN_6567;
  wire [23:0] _T_58679;
  wire [23:0] _GEN_6568;
  wire [23:0] _T_58683;
  wire [31:0] _GEN_6569;
  wire [31:0] _T_58719;
  wire [31:0] _GEN_6570;
  wire [31:0] _T_58723;
  wire [15:0] _GEN_6571;
  wire [15:0] _T_58799;
  wire [15:0] _GEN_6572;
  wire [15:0] _T_58803;
  wire [23:0] _GEN_6573;
  wire [23:0] _T_58839;
  wire [23:0] _GEN_6574;
  wire [23:0] _T_58843;
  wire [31:0] _GEN_6575;
  wire [31:0] _T_58879;
  wire [31:0] _GEN_6576;
  wire [31:0] _T_58883;
  wire [15:0] _GEN_6577;
  wire [15:0] _T_58959;
  wire [15:0] _GEN_6578;
  wire [15:0] _T_58963;
  wire [23:0] _GEN_6579;
  wire [23:0] _T_58999;
  wire [23:0] _GEN_6580;
  wire [23:0] _T_59003;
  wire [31:0] _GEN_6581;
  wire [31:0] _T_59039;
  wire [31:0] _GEN_6582;
  wire [31:0] _T_59043;
  wire [15:0] _GEN_6583;
  wire [15:0] _T_59119;
  wire [15:0] _GEN_6584;
  wire [15:0] _T_59123;
  wire [23:0] _GEN_6585;
  wire [23:0] _T_59159;
  wire [23:0] _GEN_6586;
  wire [23:0] _T_59163;
  wire [31:0] _GEN_6587;
  wire [31:0] _T_59199;
  wire [31:0] _GEN_6588;
  wire [31:0] _T_59203;
  wire [15:0] _GEN_6589;
  wire [15:0] _T_59279;
  wire [15:0] _GEN_6590;
  wire [15:0] _T_59283;
  wire [23:0] _GEN_6591;
  wire [23:0] _T_59319;
  wire [23:0] _GEN_6592;
  wire [23:0] _T_59323;
  wire [31:0] _GEN_6593;
  wire [31:0] _T_59359;
  wire [31:0] _GEN_6594;
  wire [31:0] _T_59363;
  wire [15:0] _GEN_6595;
  wire [15:0] _T_59439;
  wire [15:0] _GEN_6596;
  wire [15:0] _T_59443;
  wire [23:0] _GEN_6597;
  wire [23:0] _T_59479;
  wire [23:0] _GEN_6598;
  wire [23:0] _T_59483;
  wire [31:0] _GEN_6599;
  wire [31:0] _T_59519;
  wire [31:0] _GEN_6600;
  wire [31:0] _T_59523;
  wire [15:0] _GEN_6601;
  wire [15:0] _T_59599;
  wire [15:0] _GEN_6602;
  wire [15:0] _T_59603;
  wire [23:0] _GEN_6603;
  wire [23:0] _T_59639;
  wire [23:0] _GEN_6604;
  wire [23:0] _T_59643;
  wire [31:0] _GEN_6605;
  wire [31:0] _T_59679;
  wire [31:0] _GEN_6606;
  wire [31:0] _T_59683;
  wire [15:0] _GEN_6607;
  wire [15:0] _T_59759;
  wire [15:0] _GEN_6608;
  wire [15:0] _T_59763;
  wire [23:0] _GEN_6609;
  wire [23:0] _T_59799;
  wire [23:0] _GEN_6610;
  wire [23:0] _T_59803;
  wire [31:0] _GEN_6611;
  wire [31:0] _T_59839;
  wire [31:0] _GEN_6612;
  wire [31:0] _T_59843;
  wire [15:0] _GEN_6613;
  wire [15:0] _T_59919;
  wire [15:0] _GEN_6614;
  wire [15:0] _T_59923;
  wire [23:0] _GEN_6615;
  wire [23:0] _T_59959;
  wire [23:0] _GEN_6616;
  wire [23:0] _T_59963;
  wire [31:0] _GEN_6617;
  wire [31:0] _T_59999;
  wire [31:0] _GEN_6618;
  wire [31:0] _T_60003;
  wire [15:0] _GEN_6619;
  wire [15:0] _T_60079;
  wire [15:0] _GEN_6620;
  wire [15:0] _T_60083;
  wire [23:0] _GEN_6621;
  wire [23:0] _T_60119;
  wire [23:0] _GEN_6622;
  wire [23:0] _T_60123;
  wire [31:0] _GEN_6623;
  wire [31:0] _T_60159;
  wire [31:0] _GEN_6624;
  wire [31:0] _T_60163;
  wire [15:0] _GEN_6625;
  wire [15:0] _T_60239;
  wire [15:0] _GEN_6626;
  wire [15:0] _T_60243;
  wire [23:0] _GEN_6627;
  wire [23:0] _T_60279;
  wire [23:0] _GEN_6628;
  wire [23:0] _T_60283;
  wire [31:0] _GEN_6629;
  wire [31:0] _T_60319;
  wire [31:0] _GEN_6630;
  wire [31:0] _T_60323;
  wire  _T_60343;
  wire [7:0] _GEN_2469;
  wire  _T_60383;
  wire [7:0] _GEN_2470;
  wire  _T_60423;
  wire [7:0] _GEN_2471;
  wire  _T_60463;
  wire [7:0] _GEN_2472;
  wire [15:0] _GEN_6637;
  wire [15:0] _T_60559;
  wire [15:0] _GEN_6638;
  wire [15:0] _T_60563;
  wire [23:0] _GEN_6639;
  wire [23:0] _T_60599;
  wire [23:0] _GEN_6640;
  wire [23:0] _T_60603;
  wire [31:0] _GEN_6641;
  wire [31:0] _T_60639;
  wire [31:0] _GEN_6642;
  wire [31:0] _T_60643;
  wire [15:0] _GEN_6643;
  wire [15:0] _T_60719;
  wire [15:0] _GEN_6644;
  wire [15:0] _T_60723;
  wire [23:0] _GEN_6645;
  wire [23:0] _T_60759;
  wire [23:0] _GEN_6646;
  wire [23:0] _T_60763;
  wire [31:0] _GEN_6647;
  wire [31:0] _T_60799;
  wire [31:0] _GEN_6648;
  wire [31:0] _T_60803;
  wire [15:0] _GEN_6649;
  wire [15:0] _T_60879;
  wire [15:0] _GEN_6650;
  wire [15:0] _T_60883;
  wire [23:0] _GEN_6651;
  wire [23:0] _T_60919;
  wire [23:0] _GEN_6652;
  wire [23:0] _T_60923;
  wire [31:0] _GEN_6653;
  wire [31:0] _T_60959;
  wire [31:0] _GEN_6654;
  wire [31:0] _T_60963;
  wire [15:0] _GEN_6655;
  wire [15:0] _T_61039;
  wire [15:0] _GEN_6656;
  wire [15:0] _T_61043;
  wire [23:0] _GEN_6657;
  wire [23:0] _T_61079;
  wire [23:0] _GEN_6658;
  wire [23:0] _T_61083;
  wire [31:0] _GEN_6659;
  wire [31:0] _T_61119;
  wire [31:0] _GEN_6660;
  wire [31:0] _T_61123;
  wire [15:0] _GEN_6661;
  wire [15:0] _T_61199;
  wire [15:0] _GEN_6662;
  wire [15:0] _T_61203;
  wire [23:0] _GEN_6663;
  wire [23:0] _T_61239;
  wire [23:0] _GEN_6664;
  wire [23:0] _T_61243;
  wire [31:0] _GEN_6665;
  wire [31:0] _T_61279;
  wire [31:0] _GEN_6666;
  wire [31:0] _T_61283;
  wire [15:0] _GEN_6667;
  wire [15:0] _T_61359;
  wire [15:0] _GEN_6668;
  wire [15:0] _T_61363;
  wire [23:0] _GEN_6669;
  wire [23:0] _T_61399;
  wire [23:0] _GEN_6670;
  wire [23:0] _T_61403;
  wire [31:0] _GEN_6671;
  wire [31:0] _T_61439;
  wire [31:0] _GEN_6672;
  wire [31:0] _T_61443;
  wire [15:0] _GEN_6673;
  wire [15:0] _T_61519;
  wire [15:0] _GEN_6674;
  wire [15:0] _T_61523;
  wire [23:0] _GEN_6675;
  wire [23:0] _T_61559;
  wire [23:0] _GEN_6676;
  wire [23:0] _T_61563;
  wire [31:0] _GEN_6677;
  wire [31:0] _T_61599;
  wire [31:0] _GEN_6678;
  wire [31:0] _T_61603;
  wire [15:0] _GEN_6679;
  wire [15:0] _T_61679;
  wire [15:0] _GEN_6680;
  wire [15:0] _T_61683;
  wire [23:0] _GEN_6681;
  wire [23:0] _T_61719;
  wire [23:0] _GEN_6682;
  wire [23:0] _T_61723;
  wire [31:0] _GEN_6683;
  wire [31:0] _T_61759;
  wire [31:0] _GEN_6684;
  wire [31:0] _T_61763;
  wire [15:0] _GEN_6685;
  wire [15:0] _T_61839;
  wire [15:0] _GEN_6686;
  wire [15:0] _T_61843;
  wire [23:0] _GEN_6687;
  wire [23:0] _T_61879;
  wire [23:0] _GEN_6688;
  wire [23:0] _T_61883;
  wire [31:0] _GEN_6689;
  wire [31:0] _T_61919;
  wire [31:0] _GEN_6690;
  wire [31:0] _T_61923;
  wire [15:0] _GEN_6691;
  wire [15:0] _T_61999;
  wire [15:0] _GEN_6692;
  wire [15:0] _T_62003;
  wire [23:0] _GEN_6693;
  wire [23:0] _T_62039;
  wire [23:0] _GEN_6694;
  wire [23:0] _T_62043;
  wire [31:0] _GEN_6695;
  wire [31:0] _T_62079;
  wire [31:0] _GEN_6696;
  wire [31:0] _T_62083;
  wire  _T_62103;
  wire [7:0] _GEN_2473;
  wire  _T_62143;
  wire [7:0] _GEN_2474;
  wire  _T_62183;
  wire [7:0] _GEN_2475;
  wire  _T_62223;
  wire [7:0] _GEN_2476;
  wire [15:0] _GEN_6703;
  wire [15:0] _T_62319;
  wire [15:0] _GEN_6704;
  wire [15:0] _T_62323;
  wire [23:0] _GEN_6705;
  wire [23:0] _T_62359;
  wire [23:0] _GEN_6706;
  wire [23:0] _T_62363;
  wire [31:0] _GEN_6707;
  wire [31:0] _T_62399;
  wire [31:0] _GEN_6708;
  wire [31:0] _T_62403;
  wire [15:0] _GEN_6709;
  wire [15:0] _T_62479;
  wire [15:0] _GEN_6710;
  wire [15:0] _T_62483;
  wire [23:0] _GEN_6711;
  wire [23:0] _T_62519;
  wire [23:0] _GEN_6712;
  wire [23:0] _T_62523;
  wire [31:0] _GEN_6713;
  wire [31:0] _T_62559;
  wire [31:0] _GEN_6714;
  wire [31:0] _T_62563;
  wire [15:0] _GEN_6715;
  wire [15:0] _T_62639;
  wire [15:0] _GEN_6716;
  wire [15:0] _T_62643;
  wire [23:0] _GEN_6717;
  wire [23:0] _T_62679;
  wire [23:0] _GEN_6718;
  wire [23:0] _T_62683;
  wire [31:0] _GEN_6719;
  wire [31:0] _T_62719;
  wire [31:0] _GEN_6720;
  wire [31:0] _T_62723;
  wire [15:0] _GEN_6721;
  wire [15:0] _T_62799;
  wire [15:0] _GEN_6722;
  wire [15:0] _T_62803;
  wire [23:0] _GEN_6723;
  wire [23:0] _T_62839;
  wire [23:0] _GEN_6724;
  wire [23:0] _T_62843;
  wire [31:0] _GEN_6725;
  wire [31:0] _T_62879;
  wire [31:0] _GEN_6726;
  wire [31:0] _T_62883;
  wire [15:0] _GEN_6727;
  wire [15:0] _T_62959;
  wire [15:0] _GEN_6728;
  wire [15:0] _T_62963;
  wire [23:0] _GEN_6729;
  wire [23:0] _T_62999;
  wire [23:0] _GEN_6730;
  wire [23:0] _T_63003;
  wire [31:0] _GEN_6731;
  wire [31:0] _T_63039;
  wire [31:0] _GEN_6732;
  wire [31:0] _T_63043;
  wire [15:0] _GEN_6733;
  wire [15:0] _T_63279;
  wire [15:0] _GEN_6734;
  wire [15:0] _T_63283;
  wire [23:0] _GEN_6735;
  wire [23:0] _T_63319;
  wire [23:0] _GEN_6736;
  wire [23:0] _T_63323;
  wire [31:0] _GEN_6737;
  wire [31:0] _T_63359;
  wire [31:0] _GEN_6738;
  wire [31:0] _T_63363;
  wire  _T_63383;
  wire [7:0] _GEN_2477;
  wire  _T_63423;
  wire [7:0] _GEN_2478;
  wire  _T_63463;
  wire [7:0] _GEN_2479;
  wire  _T_63503;
  wire [7:0] _GEN_2480;
  wire [15:0] _GEN_6745;
  wire [15:0] _T_63599;
  wire [15:0] _GEN_6746;
  wire [15:0] _T_63603;
  wire [23:0] _GEN_6747;
  wire [23:0] _T_63639;
  wire [23:0] _GEN_6748;
  wire [23:0] _T_63643;
  wire [31:0] _GEN_6749;
  wire [31:0] _T_63679;
  wire [31:0] _GEN_6750;
  wire [31:0] _T_63683;
  wire  _T_63863;
  wire [9:0] _T_63864;
  wire [15:0] _GEN_6751;
  wire [15:0] _T_63959;
  wire [15:0] _GEN_6752;
  wire [15:0] _T_63963;
  wire [23:0] _GEN_6753;
  wire [23:0] _T_63999;
  wire [23:0] _GEN_6754;
  wire [23:0] _T_64003;
  wire [31:0] _GEN_6755;
  wire [31:0] _T_64039;
  wire [31:0] _GEN_6756;
  wire [31:0] _T_64043;
  wire [15:0] _GEN_6757;
  wire [15:0] _T_64119;
  wire [15:0] _GEN_6758;
  wire [15:0] _T_64123;
  wire [23:0] _GEN_6759;
  wire [23:0] _T_64159;
  wire [23:0] _GEN_6760;
  wire [23:0] _T_64163;
  wire [31:0] _GEN_6761;
  wire [31:0] _T_64199;
  wire [31:0] _GEN_6762;
  wire [31:0] _T_64203;
  wire [15:0] _GEN_6763;
  wire [15:0] _T_64439;
  wire [15:0] _GEN_6764;
  wire [15:0] _T_64443;
  wire [23:0] _GEN_6765;
  wire [23:0] _T_64479;
  wire [23:0] _GEN_6766;
  wire [23:0] _T_64483;
  wire [31:0] _GEN_6767;
  wire [31:0] _T_64519;
  wire [31:0] _GEN_6768;
  wire [31:0] _T_64523;
  wire [15:0] _GEN_6769;
  wire [15:0] _T_64599;
  wire [15:0] _GEN_6770;
  wire [15:0] _T_64603;
  wire [23:0] _GEN_6771;
  wire [23:0] _T_64639;
  wire [23:0] _GEN_6772;
  wire [23:0] _T_64643;
  wire [31:0] _GEN_6773;
  wire [31:0] _T_64679;
  wire [31:0] _GEN_6774;
  wire [31:0] _T_64683;
  wire [15:0] _GEN_6775;
  wire [15:0] _T_64759;
  wire [15:0] _GEN_6776;
  wire [15:0] _T_64763;
  wire [23:0] _GEN_6777;
  wire [23:0] _T_64799;
  wire [23:0] _GEN_6778;
  wire [23:0] _T_64803;
  wire [31:0] _GEN_6779;
  wire [31:0] _T_64839;
  wire [31:0] _GEN_6780;
  wire [31:0] _T_64843;
  wire  _T_64863;
  wire [7:0] _GEN_2482;
  wire  _T_64903;
  wire [7:0] _GEN_2483;
  wire  _T_64943;
  wire [7:0] _GEN_2484;
  wire  _T_64983;
  wire [7:0] _GEN_2485;
  wire [15:0] _GEN_6787;
  wire [15:0] _T_65079;
  wire [15:0] _GEN_6788;
  wire [15:0] _T_65083;
  wire [23:0] _GEN_6789;
  wire [23:0] _T_65119;
  wire [23:0] _GEN_6790;
  wire [23:0] _T_65123;
  wire [31:0] _GEN_6791;
  wire [31:0] _T_65159;
  wire [31:0] _GEN_6792;
  wire [31:0] _T_65163;
  wire [15:0] _GEN_6793;
  wire [15:0] _T_65239;
  wire [15:0] _GEN_6794;
  wire [15:0] _T_65243;
  wire [23:0] _GEN_6795;
  wire [23:0] _T_65279;
  wire [23:0] _GEN_6796;
  wire [23:0] _T_65283;
  wire [31:0] _GEN_6797;
  wire [31:0] _T_65319;
  wire [31:0] _GEN_6798;
  wire [31:0] _T_65323;
  wire [15:0] _GEN_6799;
  wire [15:0] _T_65399;
  wire [15:0] _GEN_6800;
  wire [15:0] _T_65403;
  wire [23:0] _GEN_6801;
  wire [23:0] _T_65439;
  wire [23:0] _GEN_6802;
  wire [23:0] _T_65443;
  wire [31:0] _GEN_6803;
  wire [31:0] _T_65479;
  wire [31:0] _GEN_6804;
  wire [31:0] _T_65483;
  wire [15:0] _GEN_6805;
  wire [15:0] _T_65559;
  wire [15:0] _GEN_6806;
  wire [15:0] _T_65563;
  wire [23:0] _GEN_6807;
  wire [23:0] _T_65599;
  wire [23:0] _GEN_6808;
  wire [23:0] _T_65603;
  wire [31:0] _GEN_6809;
  wire [31:0] _T_65639;
  wire [31:0] _GEN_6810;
  wire [31:0] _T_65643;
  wire [15:0] _GEN_6811;
  wire [15:0] _T_65719;
  wire [15:0] _GEN_6812;
  wire [15:0] _T_65723;
  wire [23:0] _GEN_6813;
  wire [23:0] _T_65759;
  wire [23:0] _GEN_6814;
  wire [23:0] _T_65763;
  wire [31:0] _GEN_6815;
  wire [31:0] _T_65799;
  wire [31:0] _GEN_6816;
  wire [31:0] _T_65803;
  wire [15:0] _GEN_6817;
  wire [15:0] _T_65879;
  wire [15:0] _GEN_6818;
  wire [15:0] _T_65883;
  wire [23:0] _GEN_6819;
  wire [23:0] _T_65919;
  wire [23:0] _GEN_6820;
  wire [23:0] _T_65923;
  wire [31:0] _GEN_6821;
  wire [31:0] _T_65959;
  wire [31:0] _GEN_6822;
  wire [31:0] _T_65963;
  wire [15:0] _GEN_6823;
  wire [15:0] _T_66039;
  wire [15:0] _GEN_6824;
  wire [15:0] _T_66043;
  wire [23:0] _GEN_6825;
  wire [23:0] _T_66079;
  wire [23:0] _GEN_6826;
  wire [23:0] _T_66083;
  wire [31:0] _GEN_6827;
  wire [31:0] _T_66119;
  wire [31:0] _GEN_6828;
  wire [31:0] _T_66123;
  wire [15:0] _GEN_6829;
  wire [15:0] _T_66199;
  wire [15:0] _GEN_6830;
  wire [15:0] _T_66203;
  wire [23:0] _GEN_6831;
  wire [23:0] _T_66239;
  wire [23:0] _GEN_6832;
  wire [23:0] _T_66243;
  wire [31:0] _GEN_6833;
  wire [31:0] _T_66279;
  wire [31:0] _GEN_6834;
  wire [31:0] _T_66283;
  wire [15:0] _GEN_6835;
  wire [15:0] _T_66359;
  wire [15:0] _GEN_6836;
  wire [15:0] _T_66363;
  wire [23:0] _GEN_6837;
  wire [23:0] _T_66399;
  wire [23:0] _GEN_6838;
  wire [23:0] _T_66403;
  wire [31:0] _GEN_6839;
  wire [31:0] _T_66439;
  wire [31:0] _GEN_6840;
  wire [31:0] _T_66443;
  wire [15:0] _GEN_6841;
  wire [15:0] _T_66519;
  wire [15:0] _GEN_6842;
  wire [15:0] _T_66523;
  wire [23:0] _GEN_6843;
  wire [23:0] _T_66559;
  wire [23:0] _GEN_6844;
  wire [23:0] _T_66563;
  wire [31:0] _GEN_6845;
  wire [31:0] _T_66599;
  wire [31:0] _GEN_6846;
  wire [31:0] _T_66603;
  wire [15:0] _GEN_6847;
  wire [15:0] _T_66839;
  wire [15:0] _GEN_6848;
  wire [15:0] _T_66843;
  wire [23:0] _GEN_6849;
  wire [23:0] _T_66879;
  wire [23:0] _GEN_6850;
  wire [23:0] _T_66883;
  wire [31:0] _GEN_6851;
  wire [31:0] _T_66919;
  wire [31:0] _GEN_6852;
  wire [31:0] _T_66923;
  wire  _T_66943;
  wire [7:0] _GEN_2486;
  wire  _T_66983;
  wire [7:0] _GEN_2487;
  wire  _T_67023;
  wire [7:0] _GEN_2488;
  wire  _T_67063;
  wire [7:0] _GEN_2489;
  wire [15:0] _GEN_6859;
  wire [15:0] _T_67159;
  wire [15:0] _GEN_6860;
  wire [15:0] _T_67163;
  wire [23:0] _GEN_6861;
  wire [23:0] _T_67199;
  wire [23:0] _GEN_6862;
  wire [23:0] _T_67203;
  wire [31:0] _GEN_6863;
  wire [31:0] _T_67239;
  wire [31:0] _GEN_6864;
  wire [31:0] _T_67243;
  wire [15:0] _GEN_6865;
  wire [15:0] _T_67479;
  wire [15:0] _GEN_6866;
  wire [15:0] _T_67483;
  wire [23:0] _GEN_6867;
  wire [23:0] _T_67519;
  wire [23:0] _GEN_6868;
  wire [23:0] _T_67523;
  wire [31:0] _GEN_6869;
  wire [31:0] _T_67559;
  wire [31:0] _GEN_6870;
  wire [31:0] _T_67563;
  wire [15:0] _GEN_6871;
  wire [15:0] _T_67639;
  wire [15:0] _GEN_6872;
  wire [15:0] _T_67643;
  wire [23:0] _GEN_6873;
  wire [23:0] _T_67679;
  wire [23:0] _GEN_6874;
  wire [23:0] _T_67683;
  wire [31:0] _GEN_6875;
  wire [31:0] _T_67719;
  wire [31:0] _GEN_6876;
  wire [31:0] _T_67723;
  wire [15:0] _GEN_6877;
  wire [15:0] _T_67799;
  wire [15:0] _GEN_6878;
  wire [15:0] _T_67803;
  wire [23:0] _GEN_6879;
  wire [23:0] _T_67839;
  wire [23:0] _GEN_6880;
  wire [23:0] _T_67843;
  wire [31:0] _GEN_6881;
  wire [31:0] _T_67879;
  wire [31:0] _GEN_6882;
  wire [31:0] _T_67883;
  wire [15:0] _GEN_6883;
  wire [15:0] _T_68119;
  wire [15:0] _GEN_6884;
  wire [15:0] _T_68123;
  wire [23:0] _GEN_6885;
  wire [23:0] _T_68159;
  wire [23:0] _GEN_6886;
  wire [23:0] _T_68163;
  wire [31:0] _GEN_6887;
  wire [31:0] _T_68199;
  wire [31:0] _GEN_6888;
  wire [31:0] _T_68203;
  wire [15:0] _GEN_6889;
  wire [15:0] _T_68279;
  wire [15:0] _GEN_6890;
  wire [15:0] _T_68283;
  wire [23:0] _GEN_6891;
  wire [23:0] _T_68319;
  wire [23:0] _GEN_6892;
  wire [23:0] _T_68323;
  wire [31:0] _GEN_6893;
  wire [31:0] _T_68359;
  wire [31:0] _GEN_6894;
  wire [31:0] _T_68363;
  wire [15:0] _GEN_6895;
  wire [15:0] _T_68439;
  wire [15:0] _GEN_6896;
  wire [15:0] _T_68443;
  wire [23:0] _GEN_6897;
  wire [23:0] _T_68479;
  wire [23:0] _GEN_6898;
  wire [23:0] _T_68483;
  wire [31:0] _GEN_6899;
  wire [31:0] _T_68519;
  wire [31:0] _GEN_6900;
  wire [31:0] _T_68523;
  wire [15:0] _GEN_6901;
  wire [15:0] _T_68599;
  wire [15:0] _GEN_6902;
  wire [15:0] _T_68603;
  wire [23:0] _GEN_6903;
  wire [23:0] _T_68639;
  wire [23:0] _GEN_6904;
  wire [23:0] _T_68643;
  wire [31:0] _GEN_6905;
  wire [31:0] _T_68679;
  wire [31:0] _GEN_6906;
  wire [31:0] _T_68683;
  wire [15:0] _GEN_6907;
  wire [15:0] _T_68759;
  wire [15:0] _GEN_6908;
  wire [15:0] _T_68763;
  wire [23:0] _GEN_6909;
  wire [23:0] _T_68799;
  wire [23:0] _GEN_6910;
  wire [23:0] _T_68803;
  wire [31:0] _GEN_6911;
  wire [31:0] _T_68839;
  wire [31:0] _GEN_6912;
  wire [31:0] _T_68843;
  wire [15:0] _GEN_6913;
  wire [15:0] _T_68919;
  wire [15:0] _GEN_6914;
  wire [15:0] _T_68923;
  wire [23:0] _GEN_6915;
  wire [23:0] _T_68959;
  wire [23:0] _GEN_6916;
  wire [23:0] _T_68963;
  wire [31:0] _GEN_6917;
  wire [31:0] _T_68999;
  wire [31:0] _GEN_6918;
  wire [31:0] _T_69003;
  wire [15:0] _GEN_6919;
  wire [15:0] _T_69079;
  wire [15:0] _GEN_6920;
  wire [15:0] _T_69083;
  wire [23:0] _GEN_6921;
  wire [23:0] _T_69119;
  wire [23:0] _GEN_6922;
  wire [23:0] _T_69123;
  wire [31:0] _GEN_6923;
  wire [31:0] _T_69159;
  wire [31:0] _GEN_6924;
  wire [31:0] _T_69163;
  wire  _T_69183;
  wire [15:0] _GEN_6925;
  wire [15:0] _T_69279;
  wire [15:0] _GEN_6926;
  wire [15:0] _T_69283;
  wire [23:0] _GEN_6927;
  wire [23:0] _T_69319;
  wire [23:0] _GEN_6928;
  wire [23:0] _T_69323;
  wire [31:0] _GEN_6929;
  wire [31:0] _T_69359;
  wire [31:0] _GEN_6930;
  wire [31:0] _T_69363;
  wire [15:0] _GEN_6931;
  wire [15:0] _T_69439;
  wire [15:0] _GEN_6932;
  wire [15:0] _T_69443;
  wire [23:0] _GEN_6933;
  wire [23:0] _T_69479;
  wire [23:0] _GEN_6934;
  wire [23:0] _T_69483;
  wire [31:0] _GEN_6935;
  wire [31:0] _T_69519;
  wire [31:0] _GEN_6936;
  wire [31:0] _T_69523;
  wire [15:0] _GEN_6937;
  wire [15:0] _T_69599;
  wire [15:0] _GEN_6938;
  wire [15:0] _T_69603;
  wire [23:0] _GEN_6939;
  wire [23:0] _T_69639;
  wire [23:0] _GEN_6940;
  wire [23:0] _T_69643;
  wire [31:0] _GEN_6941;
  wire [31:0] _T_69679;
  wire [31:0] _GEN_6942;
  wire [31:0] _T_69683;
  wire [15:0] _GEN_6943;
  wire [15:0] _T_69759;
  wire [15:0] _GEN_6944;
  wire [15:0] _T_69763;
  wire [23:0] _GEN_6945;
  wire [23:0] _T_69799;
  wire [23:0] _GEN_6946;
  wire [23:0] _T_69803;
  wire [31:0] _GEN_6947;
  wire [31:0] _T_69839;
  wire [31:0] _GEN_6948;
  wire [31:0] _T_69843;
  wire [15:0] _GEN_6949;
  wire [15:0] _T_69919;
  wire [15:0] _GEN_6950;
  wire [15:0] _T_69923;
  wire [23:0] _GEN_6951;
  wire [23:0] _T_69959;
  wire [23:0] _GEN_6952;
  wire [23:0] _T_69963;
  wire [31:0] _GEN_6953;
  wire [31:0] _T_69999;
  wire [31:0] _GEN_6954;
  wire [31:0] _T_70003;
  wire [15:0] _GEN_6955;
  wire [15:0] _T_70079;
  wire [15:0] _GEN_6956;
  wire [15:0] _T_70083;
  wire [23:0] _GEN_6957;
  wire [23:0] _T_70119;
  wire [23:0] _GEN_6958;
  wire [23:0] _T_70123;
  wire [31:0] _GEN_6959;
  wire [31:0] _T_70159;
  wire [31:0] _GEN_6960;
  wire [31:0] _T_70163;
  wire [15:0] _GEN_6961;
  wire [15:0] _T_70239;
  wire [15:0] _GEN_6962;
  wire [15:0] _T_70243;
  wire [23:0] _GEN_6963;
  wire [23:0] _T_70279;
  wire [23:0] _GEN_6964;
  wire [23:0] _T_70283;
  wire [31:0] _GEN_6965;
  wire [31:0] _T_70319;
  wire [31:0] _GEN_6966;
  wire [31:0] _T_70323;
  wire [15:0] _GEN_6967;
  wire [15:0] _T_70399;
  wire [15:0] _GEN_6968;
  wire [15:0] _T_70403;
  wire [23:0] _GEN_6969;
  wire [23:0] _T_70439;
  wire [23:0] _GEN_6970;
  wire [23:0] _T_70443;
  wire [31:0] _GEN_6971;
  wire [31:0] _T_70479;
  wire [31:0] _GEN_6972;
  wire [31:0] _T_70483;
  wire [15:0] _GEN_6973;
  wire [15:0] _T_70559;
  wire [15:0] _GEN_6974;
  wire [15:0] _T_70563;
  wire [23:0] _GEN_6975;
  wire [23:0] _T_70599;
  wire [23:0] _GEN_6976;
  wire [23:0] _T_70603;
  wire [31:0] _GEN_6977;
  wire [31:0] _T_70639;
  wire [31:0] _GEN_6978;
  wire [31:0] _T_70643;
  wire [15:0] _GEN_6979;
  wire [15:0] _T_70719;
  wire [15:0] _GEN_6980;
  wire [15:0] _T_70723;
  wire [23:0] _GEN_6981;
  wire [23:0] _T_70759;
  wire [23:0] _GEN_6982;
  wire [23:0] _T_70763;
  wire [31:0] _GEN_6983;
  wire [31:0] _T_70799;
  wire [31:0] _GEN_6984;
  wire [31:0] _T_70803;
  wire [15:0] _GEN_6985;
  wire [15:0] _T_70879;
  wire [15:0] _GEN_6986;
  wire [15:0] _T_70883;
  wire [23:0] _GEN_6987;
  wire [23:0] _T_70919;
  wire [23:0] _GEN_6988;
  wire [23:0] _T_70923;
  wire [31:0] _GEN_6989;
  wire [31:0] _T_70959;
  wire [31:0] _GEN_6990;
  wire [31:0] _T_70963;
  wire [15:0] _GEN_6991;
  wire [15:0] _T_71039;
  wire [15:0] _GEN_6992;
  wire [15:0] _T_71043;
  wire [23:0] _GEN_6993;
  wire [23:0] _T_71079;
  wire [23:0] _GEN_6994;
  wire [23:0] _T_71083;
  wire [31:0] _GEN_6995;
  wire [31:0] _T_71119;
  wire [31:0] _GEN_6996;
  wire [31:0] _T_71123;
  wire [15:0] _GEN_6997;
  wire [15:0] _T_71199;
  wire [15:0] _GEN_6998;
  wire [15:0] _T_71203;
  wire [23:0] _GEN_6999;
  wire [23:0] _T_71239;
  wire [23:0] _GEN_7000;
  wire [23:0] _T_71243;
  wire [31:0] _GEN_7001;
  wire [31:0] _T_71279;
  wire [31:0] _GEN_7002;
  wire [31:0] _T_71283;
  wire [15:0] _GEN_7003;
  wire [15:0] _T_71359;
  wire [15:0] _GEN_7004;
  wire [15:0] _T_71363;
  wire [23:0] _GEN_7005;
  wire [23:0] _T_71399;
  wire [23:0] _GEN_7006;
  wire [23:0] _T_71403;
  wire [31:0] _GEN_7007;
  wire [31:0] _T_71439;
  wire [31:0] _GEN_7008;
  wire [31:0] _T_71443;
  wire [15:0] _GEN_7009;
  wire [15:0] _T_71519;
  wire [15:0] _GEN_7010;
  wire [15:0] _T_71523;
  wire [23:0] _GEN_7011;
  wire [23:0] _T_71559;
  wire [23:0] _GEN_7012;
  wire [23:0] _T_71563;
  wire [31:0] _GEN_7013;
  wire [31:0] _T_71599;
  wire [31:0] _GEN_7014;
  wire [31:0] _T_71603;
  wire [15:0] _GEN_7015;
  wire [15:0] _T_71679;
  wire [15:0] _GEN_7016;
  wire [15:0] _T_71683;
  wire [23:0] _GEN_7017;
  wire [23:0] _T_71719;
  wire [23:0] _GEN_7018;
  wire [23:0] _T_71723;
  wire [31:0] _GEN_7019;
  wire [31:0] _T_71759;
  wire [31:0] _GEN_7020;
  wire [31:0] _T_71763;
  wire [15:0] _GEN_7021;
  wire [15:0] _T_71839;
  wire [15:0] _GEN_7022;
  wire [15:0] _T_71843;
  wire [23:0] _GEN_7023;
  wire [23:0] _T_71879;
  wire [23:0] _GEN_7024;
  wire [23:0] _T_71883;
  wire [31:0] _GEN_7025;
  wire [31:0] _T_71919;
  wire [31:0] _GEN_7026;
  wire [31:0] _T_71923;
  wire [15:0] _GEN_7027;
  wire [15:0] _T_72159;
  wire [15:0] _GEN_7028;
  wire [15:0] _T_72163;
  wire [23:0] _GEN_7029;
  wire [23:0] _T_72199;
  wire [23:0] _GEN_7030;
  wire [23:0] _T_72203;
  wire [31:0] _GEN_7031;
  wire [31:0] _T_72239;
  wire [31:0] _GEN_7032;
  wire [31:0] _T_72243;
  wire  _T_72263;
  wire [7:0] _GEN_2491;
  wire  _T_72303;
  wire [7:0] _GEN_2492;
  wire  _T_72343;
  wire [7:0] _GEN_2493;
  wire  _T_72383;
  wire [7:0] _GEN_2494;
  wire [15:0] _GEN_7039;
  wire [15:0] _T_72479;
  wire [15:0] _GEN_7040;
  wire [15:0] _T_72483;
  wire [23:0] _GEN_7041;
  wire [23:0] _T_72519;
  wire [23:0] _GEN_7042;
  wire [23:0] _T_72523;
  wire [31:0] _GEN_7043;
  wire [31:0] _T_72559;
  wire [31:0] _GEN_7044;
  wire [31:0] _T_72563;
  wire [15:0] _GEN_7045;
  wire [15:0] _T_72799;
  wire [15:0] _GEN_7046;
  wire [15:0] _T_72803;
  wire [23:0] _GEN_7047;
  wire [23:0] _T_72839;
  wire [23:0] _GEN_7048;
  wire [23:0] _T_72843;
  wire [31:0] _GEN_7049;
  wire [31:0] _T_72879;
  wire [31:0] _GEN_7050;
  wire [31:0] _T_72883;
  wire [15:0] _GEN_7051;
  wire [15:0] _T_72959;
  wire [15:0] _GEN_7052;
  wire [15:0] _T_72963;
  wire [23:0] _GEN_7053;
  wire [23:0] _T_72999;
  wire [23:0] _GEN_7054;
  wire [23:0] _T_73003;
  wire [31:0] _GEN_7055;
  wire [31:0] _T_73039;
  wire [31:0] _GEN_7056;
  wire [31:0] _T_73043;
  wire [15:0] _GEN_7057;
  wire [15:0] _T_73119;
  wire [15:0] _GEN_7058;
  wire [15:0] _T_73123;
  wire [23:0] _GEN_7059;
  wire [23:0] _T_73159;
  wire [23:0] _GEN_7060;
  wire [23:0] _T_73163;
  wire [31:0] _GEN_7061;
  wire [31:0] _T_73199;
  wire [31:0] _GEN_7062;
  wire [31:0] _T_73203;
  wire [15:0] _GEN_7063;
  wire [15:0] _T_73279;
  wire [15:0] _GEN_7064;
  wire [15:0] _T_73283;
  wire [23:0] _GEN_7065;
  wire [23:0] _T_73319;
  wire [23:0] _GEN_7066;
  wire [23:0] _T_73323;
  wire [31:0] _GEN_7067;
  wire [31:0] _T_73359;
  wire [31:0] _GEN_7068;
  wire [31:0] _T_73363;
  wire [15:0] _GEN_7069;
  wire [15:0] _T_73439;
  wire [15:0] _GEN_7070;
  wire [15:0] _T_73443;
  wire [23:0] _GEN_7071;
  wire [23:0] _T_73479;
  wire [23:0] _GEN_7072;
  wire [23:0] _T_73483;
  wire [31:0] _GEN_7073;
  wire [31:0] _T_73519;
  wire [31:0] _GEN_7074;
  wire [31:0] _T_73523;
  wire [15:0] _GEN_7075;
  wire [15:0] _T_73599;
  wire [15:0] _GEN_7076;
  wire [15:0] _T_73603;
  wire [23:0] _GEN_7077;
  wire [23:0] _T_73639;
  wire [23:0] _GEN_7078;
  wire [23:0] _T_73643;
  wire [31:0] _GEN_7079;
  wire [31:0] _T_73679;
  wire [31:0] _GEN_7080;
  wire [31:0] _T_73683;
  wire [15:0] _GEN_7081;
  wire [15:0] _T_73759;
  wire [15:0] _GEN_7082;
  wire [15:0] _T_73763;
  wire [23:0] _GEN_7083;
  wire [23:0] _T_73799;
  wire [23:0] _GEN_7084;
  wire [23:0] _T_73803;
  wire [31:0] _GEN_7085;
  wire [31:0] _T_73839;
  wire [31:0] _GEN_7086;
  wire [31:0] _T_73843;
  wire [15:0] _GEN_7087;
  wire [15:0] _T_73919;
  wire [15:0] _GEN_7088;
  wire [15:0] _T_73923;
  wire [23:0] _GEN_7089;
  wire [23:0] _T_73959;
  wire [23:0] _GEN_7090;
  wire [23:0] _T_73963;
  wire [31:0] _GEN_7091;
  wire [31:0] _T_73999;
  wire [31:0] _GEN_7092;
  wire [31:0] _T_74003;
  wire [15:0] _GEN_7093;
  wire [15:0] _T_74079;
  wire [15:0] _GEN_7094;
  wire [15:0] _T_74083;
  wire [23:0] _GEN_7095;
  wire [23:0] _T_74119;
  wire [23:0] _GEN_7096;
  wire [23:0] _T_74123;
  wire [31:0] _GEN_7097;
  wire [31:0] _T_74159;
  wire [31:0] _GEN_7098;
  wire [31:0] _T_74163;
  wire [15:0] _GEN_7099;
  wire [15:0] _T_74239;
  wire [15:0] _GEN_7100;
  wire [15:0] _T_74243;
  wire [23:0] _GEN_7101;
  wire [23:0] _T_74279;
  wire [23:0] _GEN_7102;
  wire [23:0] _T_74283;
  wire [31:0] _GEN_7103;
  wire [31:0] _T_74319;
  wire [31:0] _GEN_7104;
  wire [31:0] _T_74323;
  wire [15:0] _GEN_7105;
  wire [15:0] _T_74399;
  wire [15:0] _GEN_7106;
  wire [15:0] _T_74403;
  wire [23:0] _GEN_7107;
  wire [23:0] _T_74439;
  wire [23:0] _GEN_7108;
  wire [23:0] _T_74443;
  wire [31:0] _GEN_7109;
  wire [31:0] _T_74479;
  wire [31:0] _GEN_7110;
  wire [31:0] _T_74483;
  wire [15:0] _GEN_7111;
  wire [15:0] _T_74599;
  wire [15:0] _GEN_7112;
  wire [15:0] _T_74603;
  wire [23:0] _GEN_7113;
  wire [23:0] _T_74639;
  wire [23:0] _GEN_7114;
  wire [23:0] _T_74643;
  wire [31:0] _GEN_7115;
  wire [31:0] _T_74679;
  wire [31:0] _GEN_7116;
  wire [31:0] _T_74683;
  wire [15:0] _GEN_7117;
  wire [15:0] _T_74759;
  wire [15:0] _GEN_7118;
  wire [15:0] _T_74763;
  wire [23:0] _GEN_7119;
  wire [23:0] _T_74799;
  wire [23:0] _GEN_7120;
  wire [23:0] _T_74803;
  wire [31:0] _GEN_7121;
  wire [31:0] _T_74839;
  wire [31:0] _GEN_7122;
  wire [31:0] _T_74843;
  wire [15:0] _GEN_7123;
  wire [15:0] _T_74919;
  wire [15:0] _GEN_7124;
  wire [15:0] _T_74923;
  wire [23:0] _GEN_7125;
  wire [23:0] _T_74959;
  wire [23:0] _GEN_7126;
  wire [23:0] _T_74963;
  wire [31:0] _GEN_7127;
  wire [31:0] _T_74999;
  wire [31:0] _GEN_7128;
  wire [31:0] _T_75003;
  wire [15:0] _GEN_7129;
  wire [15:0] _T_75079;
  wire [15:0] _GEN_7130;
  wire [15:0] _T_75083;
  wire [23:0] _GEN_7131;
  wire [23:0] _T_75119;
  wire [23:0] _GEN_7132;
  wire [23:0] _T_75123;
  wire [31:0] _GEN_7133;
  wire [31:0] _T_75159;
  wire [31:0] _GEN_7134;
  wire [31:0] _T_75163;
  wire  _T_75183;
  wire [7:0] _GEN_2495;
  wire  _T_75223;
  wire [7:0] _GEN_2496;
  wire  _T_75263;
  wire [7:0] _GEN_2497;
  wire  _T_75303;
  wire [7:0] _GEN_2498;
  wire [15:0] _GEN_7141;
  wire [15:0] _T_75399;
  wire [15:0] _GEN_7142;
  wire [15:0] _T_75403;
  wire [23:0] _GEN_7143;
  wire [23:0] _T_75439;
  wire [23:0] _GEN_7144;
  wire [23:0] _T_75443;
  wire [31:0] _GEN_7145;
  wire [31:0] _T_75479;
  wire [31:0] _GEN_7146;
  wire [31:0] _T_75483;
  wire [15:0] _GEN_7147;
  wire [15:0] _T_75559;
  wire [15:0] _GEN_7148;
  wire [15:0] _T_75563;
  wire [23:0] _GEN_7149;
  wire [23:0] _T_75599;
  wire [23:0] _GEN_7150;
  wire [23:0] _T_75603;
  wire [31:0] _GEN_7151;
  wire [31:0] _T_75639;
  wire [31:0] _GEN_7152;
  wire [31:0] _T_75643;
  wire [15:0] _GEN_7153;
  wire [15:0] _T_75719;
  wire [15:0] _GEN_7154;
  wire [15:0] _T_75723;
  wire [23:0] _GEN_7155;
  wire [23:0] _T_75759;
  wire [23:0] _GEN_7156;
  wire [23:0] _T_75763;
  wire [31:0] _GEN_7157;
  wire [31:0] _T_75799;
  wire [31:0] _GEN_7158;
  wire [31:0] _T_75803;
  wire [15:0] _GEN_7159;
  wire [15:0] _T_75879;
  wire [15:0] _GEN_7160;
  wire [15:0] _T_75883;
  wire [23:0] _GEN_7161;
  wire [23:0] _T_75919;
  wire [23:0] _GEN_7162;
  wire [23:0] _T_75923;
  wire [31:0] _GEN_7163;
  wire [31:0] _T_75959;
  wire [31:0] _GEN_7164;
  wire [31:0] _T_75963;
  wire [15:0] _GEN_7165;
  wire [15:0] _T_76039;
  wire [15:0] _GEN_7166;
  wire [15:0] _T_76043;
  wire [23:0] _GEN_7167;
  wire [23:0] _T_76079;
  wire [23:0] _GEN_7168;
  wire [23:0] _T_76083;
  wire [31:0] _GEN_7169;
  wire [31:0] _T_76119;
  wire [31:0] _GEN_7170;
  wire [31:0] _T_76123;
  wire [15:0] _GEN_7171;
  wire [15:0] _T_76199;
  wire [15:0] _GEN_7172;
  wire [15:0] _T_76203;
  wire [23:0] _GEN_7173;
  wire [23:0] _T_76239;
  wire [23:0] _GEN_7174;
  wire [23:0] _T_76243;
  wire [31:0] _GEN_7175;
  wire [31:0] _T_76279;
  wire [31:0] _GEN_7176;
  wire [31:0] _T_76283;
  wire [15:0] _GEN_7177;
  wire [15:0] _T_76359;
  wire [15:0] _GEN_7178;
  wire [15:0] _T_76363;
  wire [23:0] _GEN_7179;
  wire [23:0] _T_76399;
  wire [23:0] _GEN_7180;
  wire [23:0] _T_76403;
  wire [31:0] _GEN_7181;
  wire [31:0] _T_76439;
  wire [31:0] _GEN_7182;
  wire [31:0] _T_76443;
  wire [15:0] _GEN_7183;
  wire [15:0] _T_76519;
  wire [15:0] _GEN_7184;
  wire [15:0] _T_76523;
  wire [23:0] _GEN_7185;
  wire [23:0] _T_76559;
  wire [23:0] _GEN_7186;
  wire [23:0] _T_76563;
  wire [31:0] _GEN_7187;
  wire [31:0] _T_76599;
  wire [31:0] _GEN_7188;
  wire [31:0] _T_76603;
  wire [15:0] _GEN_7189;
  wire [15:0] _T_76679;
  wire [15:0] _GEN_7190;
  wire [15:0] _T_76683;
  wire [23:0] _GEN_7191;
  wire [23:0] _T_76719;
  wire [23:0] _GEN_7192;
  wire [23:0] _T_76723;
  wire [31:0] _GEN_7193;
  wire [31:0] _T_76759;
  wire [31:0] _GEN_7194;
  wire [31:0] _T_76763;
  wire [15:0] _GEN_7195;
  wire [15:0] _T_76839;
  wire [15:0] _GEN_7196;
  wire [15:0] _T_76843;
  wire [23:0] _GEN_7197;
  wire [23:0] _T_76879;
  wire [23:0] _GEN_7198;
  wire [23:0] _T_76883;
  wire [31:0] _GEN_7199;
  wire [31:0] _T_76919;
  wire [31:0] _GEN_7200;
  wire [31:0] _T_76923;
  wire [15:0] _GEN_7201;
  wire [15:0] _T_76999;
  wire [15:0] _GEN_7202;
  wire [15:0] _T_77003;
  wire [23:0] _GEN_7203;
  wire [23:0] _T_77039;
  wire [23:0] _GEN_7204;
  wire [23:0] _T_77043;
  wire [31:0] _GEN_7205;
  wire [31:0] _T_77079;
  wire [31:0] _GEN_7206;
  wire [31:0] _T_77083;
  wire [15:0] _GEN_7207;
  wire [15:0] _T_77159;
  wire [15:0] _GEN_7208;
  wire [15:0] _T_77163;
  wire [23:0] _GEN_7209;
  wire [23:0] _T_77199;
  wire [23:0] _GEN_7210;
  wire [23:0] _T_77203;
  wire [31:0] _GEN_7211;
  wire [31:0] _T_77239;
  wire [31:0] _GEN_7212;
  wire [31:0] _T_77243;
  wire  _T_77263;
  wire [7:0] _GEN_2499;
  wire  _T_77303;
  wire [7:0] _GEN_2500;
  wire  _T_77343;
  wire [7:0] _GEN_2501;
  wire  _T_77383;
  wire [7:0] _GEN_2502;
  wire [15:0] _GEN_7219;
  wire [15:0] _T_77479;
  wire [15:0] _GEN_7220;
  wire [15:0] _T_77483;
  wire [23:0] _GEN_7221;
  wire [23:0] _T_77519;
  wire [23:0] _GEN_7222;
  wire [23:0] _T_77523;
  wire [31:0] _GEN_7223;
  wire [31:0] _T_77559;
  wire [31:0] _GEN_7224;
  wire [31:0] _T_77563;
  wire [15:0] _GEN_7225;
  wire [15:0] _T_77639;
  wire [15:0] _GEN_7226;
  wire [15:0] _T_77643;
  wire [23:0] _GEN_7227;
  wire [23:0] _T_77679;
  wire [23:0] _GEN_7228;
  wire [23:0] _T_77683;
  wire [31:0] _GEN_7229;
  wire [31:0] _T_77719;
  wire [31:0] _GEN_7230;
  wire [31:0] _T_77723;
  wire [15:0] _GEN_7231;
  wire [15:0] _T_77799;
  wire [15:0] _GEN_7232;
  wire [15:0] _T_77803;
  wire [23:0] _GEN_7233;
  wire [23:0] _T_77839;
  wire [23:0] _GEN_7234;
  wire [23:0] _T_77843;
  wire [31:0] _GEN_7235;
  wire [31:0] _T_77879;
  wire [31:0] _GEN_7236;
  wire [31:0] _T_77883;
  wire [15:0] _GEN_7237;
  wire [15:0] _T_77959;
  wire [15:0] _GEN_7238;
  wire [15:0] _T_77963;
  wire [23:0] _GEN_7239;
  wire [23:0] _T_77999;
  wire [23:0] _GEN_7240;
  wire [23:0] _T_78003;
  wire [31:0] _GEN_7241;
  wire [31:0] _T_78039;
  wire [31:0] _GEN_7242;
  wire [31:0] _T_78043;
  wire [15:0] _GEN_7243;
  wire [15:0] _T_78119;
  wire [15:0] _GEN_7244;
  wire [15:0] _T_78123;
  wire [23:0] _GEN_7245;
  wire [23:0] _T_78159;
  wire [23:0] _GEN_7246;
  wire [23:0] _T_78163;
  wire [31:0] _GEN_7247;
  wire [31:0] _T_78199;
  wire [31:0] _GEN_7248;
  wire [31:0] _T_78203;
  wire [15:0] _GEN_7249;
  wire [15:0] _T_78279;
  wire [15:0] _GEN_7250;
  wire [15:0] _T_78283;
  wire [23:0] _GEN_7251;
  wire [23:0] _T_78319;
  wire [23:0] _GEN_7252;
  wire [23:0] _T_78323;
  wire [31:0] _GEN_7253;
  wire [31:0] _T_78359;
  wire [31:0] _GEN_7254;
  wire [31:0] _T_78363;
  wire [15:0] _GEN_7255;
  wire [15:0] _T_78439;
  wire [15:0] _GEN_7256;
  wire [15:0] _T_78443;
  wire [23:0] _GEN_7257;
  wire [23:0] _T_78479;
  wire [23:0] _GEN_7258;
  wire [23:0] _T_78483;
  wire [31:0] _GEN_7259;
  wire [31:0] _T_78519;
  wire [31:0] _GEN_7260;
  wire [31:0] _T_78523;
  wire [15:0] _GEN_7261;
  wire [15:0] _T_78599;
  wire [15:0] _GEN_7262;
  wire [15:0] _T_78603;
  wire [23:0] _GEN_7263;
  wire [23:0] _T_78639;
  wire [23:0] _GEN_7264;
  wire [23:0] _T_78643;
  wire [31:0] _GEN_7265;
  wire [31:0] _T_78679;
  wire [31:0] _GEN_7266;
  wire [31:0] _T_78683;
  wire [15:0] _GEN_7267;
  wire [15:0] _T_78759;
  wire [15:0] _GEN_7268;
  wire [15:0] _T_78763;
  wire [23:0] _GEN_7269;
  wire [23:0] _T_78799;
  wire [23:0] _GEN_7270;
  wire [23:0] _T_78803;
  wire [31:0] _GEN_7271;
  wire [31:0] _T_78839;
  wire [31:0] _GEN_7272;
  wire [31:0] _T_78843;
  wire [15:0] _GEN_7273;
  wire [15:0] _T_79079;
  wire [15:0] _GEN_7274;
  wire [15:0] _T_79083;
  wire [23:0] _GEN_7275;
  wire [23:0] _T_79119;
  wire [23:0] _GEN_7276;
  wire [23:0] _T_79123;
  wire [31:0] _GEN_7277;
  wire [31:0] _T_79159;
  wire [31:0] _GEN_7278;
  wire [31:0] _T_79163;
  wire [15:0] _GEN_7279;
  wire [15:0] _T_79239;
  wire [15:0] _GEN_7280;
  wire [15:0] _T_79243;
  wire [23:0] _GEN_7281;
  wire [23:0] _T_79279;
  wire [23:0] _GEN_7282;
  wire [23:0] _T_79283;
  wire [31:0] _GEN_7283;
  wire [31:0] _T_79319;
  wire [31:0] _GEN_7284;
  wire [31:0] _T_79323;
  wire [15:0] _GEN_7285;
  wire [15:0] _T_79399;
  wire [15:0] _GEN_7286;
  wire [15:0] _T_79403;
  wire [23:0] _GEN_7287;
  wire [23:0] _T_79439;
  wire [23:0] _GEN_7288;
  wire [23:0] _T_79443;
  wire [31:0] _GEN_7289;
  wire [31:0] _T_79479;
  wire [31:0] _GEN_7290;
  wire [31:0] _T_79483;
  wire [15:0] _GEN_7291;
  wire [15:0] _T_79559;
  wire [15:0] _GEN_7292;
  wire [15:0] _T_79563;
  wire [23:0] _GEN_7293;
  wire [23:0] _T_79599;
  wire [23:0] _GEN_7294;
  wire [23:0] _T_79603;
  wire [31:0] _GEN_7295;
  wire [31:0] _T_79639;
  wire [31:0] _GEN_7296;
  wire [31:0] _T_79643;
  wire [15:0] _GEN_7297;
  wire [15:0] _T_79719;
  wire [15:0] _GEN_7298;
  wire [15:0] _T_79723;
  wire [23:0] _GEN_7299;
  wire [23:0] _T_79759;
  wire [23:0] _GEN_7300;
  wire [23:0] _T_79763;
  wire [31:0] _GEN_7301;
  wire [31:0] _T_79799;
  wire [31:0] _GEN_7302;
  wire [31:0] _T_79803;
  wire [15:0] _GEN_7303;
  wire [15:0] _T_79879;
  wire [15:0] _GEN_7304;
  wire [15:0] _T_79883;
  wire [23:0] _GEN_7305;
  wire [23:0] _T_79919;
  wire [23:0] _GEN_7306;
  wire [23:0] _T_79923;
  wire [31:0] _GEN_7307;
  wire [31:0] _T_79959;
  wire [31:0] _GEN_7308;
  wire [31:0] _T_79963;
  wire [15:0] _GEN_7309;
  wire [15:0] _T_80199;
  wire [15:0] _GEN_7310;
  wire [15:0] _T_80203;
  wire [23:0] _GEN_7311;
  wire [23:0] _T_80239;
  wire [23:0] _GEN_7312;
  wire [23:0] _T_80243;
  wire [31:0] _GEN_7313;
  wire [31:0] _T_80279;
  wire [31:0] _GEN_7314;
  wire [31:0] _T_80283;
  wire [15:0] _GEN_7315;
  wire [15:0] _T_80359;
  wire [15:0] _GEN_7316;
  wire [15:0] _T_80363;
  wire [23:0] _GEN_7317;
  wire [23:0] _T_80399;
  wire [23:0] _GEN_7318;
  wire [23:0] _T_80403;
  wire [31:0] _GEN_7319;
  wire [31:0] _T_80439;
  wire [31:0] _GEN_7320;
  wire [31:0] _T_80443;
  wire [15:0] _GEN_7321;
  wire [15:0] _T_80519;
  wire [15:0] _GEN_7322;
  wire [15:0] _T_80523;
  wire [23:0] _GEN_7323;
  wire [23:0] _T_80559;
  wire [23:0] _GEN_7324;
  wire [23:0] _T_80563;
  wire [31:0] _GEN_7325;
  wire [31:0] _T_80599;
  wire [31:0] _GEN_7326;
  wire [31:0] _T_80603;
  wire [15:0] _GEN_7327;
  wire [15:0] _T_80679;
  wire [15:0] _GEN_7328;
  wire [15:0] _T_80683;
  wire [23:0] _GEN_7329;
  wire [23:0] _T_80719;
  wire [23:0] _GEN_7330;
  wire [23:0] _T_80723;
  wire [31:0] _GEN_7331;
  wire [31:0] _T_80759;
  wire [31:0] _GEN_7332;
  wire [31:0] _T_80763;
  wire [15:0] _GEN_7333;
  wire [15:0] _T_80839;
  wire [15:0] _GEN_7334;
  wire [15:0] _T_80843;
  wire [23:0] _GEN_7335;
  wire [23:0] _T_80879;
  wire [23:0] _GEN_7336;
  wire [23:0] _T_80883;
  wire [31:0] _GEN_7337;
  wire [31:0] _T_80919;
  wire [31:0] _GEN_7338;
  wire [31:0] _T_80923;
  wire [15:0] _GEN_7339;
  wire [15:0] _T_80999;
  wire [15:0] _GEN_7340;
  wire [15:0] _T_81003;
  wire [23:0] _GEN_7341;
  wire [23:0] _T_81039;
  wire [23:0] _GEN_7342;
  wire [23:0] _T_81043;
  wire [31:0] _GEN_7343;
  wire [31:0] _T_81079;
  wire [31:0] _GEN_7344;
  wire [31:0] _T_81083;
  wire [15:0] _GEN_7345;
  wire [15:0] _T_81159;
  wire [15:0] _GEN_7346;
  wire [15:0] _T_81163;
  wire [23:0] _GEN_7347;
  wire [23:0] _T_81199;
  wire [23:0] _GEN_7348;
  wire [23:0] _T_81203;
  wire [31:0] _GEN_7349;
  wire [31:0] _T_81239;
  wire [31:0] _GEN_7350;
  wire [31:0] _T_81243;
  wire [15:0] _GEN_7351;
  wire [15:0] _T_81319;
  wire [15:0] _GEN_7352;
  wire [15:0] _T_81323;
  wire [23:0] _GEN_7353;
  wire [23:0] _T_81359;
  wire [23:0] _GEN_7354;
  wire [23:0] _T_81363;
  wire [31:0] _GEN_7355;
  wire [31:0] _T_81399;
  wire [31:0] _GEN_7356;
  wire [31:0] _T_81403;
  wire [15:0] _GEN_7357;
  wire [15:0] _T_81479;
  wire [15:0] _GEN_7358;
  wire [15:0] _T_81483;
  wire [23:0] _GEN_7359;
  wire [23:0] _T_81519;
  wire [23:0] _GEN_7360;
  wire [23:0] _T_81523;
  wire [31:0] _GEN_7361;
  wire [31:0] _T_81559;
  wire [31:0] _GEN_7362;
  wire [31:0] _T_81563;
  wire [15:0] _GEN_7363;
  wire [15:0] _T_81639;
  wire [15:0] _GEN_7364;
  wire [15:0] _T_81643;
  wire [23:0] _GEN_7365;
  wire [23:0] _T_81679;
  wire [23:0] _GEN_7366;
  wire [23:0] _T_81683;
  wire [31:0] _GEN_7367;
  wire [31:0] _T_81719;
  wire [31:0] _GEN_7368;
  wire [31:0] _T_81723;
  wire [15:0] _GEN_7369;
  wire [15:0] _T_81799;
  wire [15:0] _GEN_7370;
  wire [15:0] _T_81803;
  wire [23:0] _GEN_7371;
  wire [23:0] _T_81839;
  wire [23:0] _GEN_7372;
  wire [23:0] _T_81843;
  wire [31:0] _GEN_7373;
  wire [31:0] _T_81879;
  wire [31:0] _GEN_7374;
  wire [31:0] _T_81883;
  wire  _T_81903;
  wire [7:0] _GEN_2503;
  wire  _T_81943;
  wire [7:0] _GEN_2504;
  wire  _T_81983;
  wire [7:0] _GEN_2505;
  wire  _T_82023;
  wire [7:0] _GEN_2506;
  wire [15:0] _GEN_7381;
  wire [15:0] _T_82119;
  wire [15:0] _GEN_7382;
  wire [15:0] _T_82123;
  wire [23:0] _GEN_7383;
  wire [23:0] _T_82159;
  wire [23:0] _GEN_7384;
  wire [23:0] _T_82163;
  wire [31:0] _GEN_7385;
  wire [31:0] _T_82199;
  wire [31:0] _GEN_7386;
  wire [31:0] _T_82203;
  wire  _T_82223;
  wire [7:0] _GEN_2507;
  wire  _T_82263;
  wire [7:0] _GEN_2508;
  wire  _T_82303;
  wire [7:0] _GEN_2509;
  wire  _T_82343;
  wire [7:0] _GEN_2510;
  wire [15:0] _GEN_7393;
  wire [15:0] _T_82439;
  wire [15:0] _GEN_7394;
  wire [15:0] _T_82443;
  wire [23:0] _GEN_7395;
  wire [23:0] _T_82479;
  wire [23:0] _GEN_7396;
  wire [23:0] _T_82483;
  wire [31:0] _GEN_7397;
  wire [31:0] _T_82519;
  wire [31:0] _GEN_7398;
  wire [31:0] _T_82523;
  wire [15:0] _GEN_7399;
  wire [15:0] _T_82599;
  wire [15:0] _GEN_7400;
  wire [15:0] _T_82603;
  wire [23:0] _GEN_7401;
  wire [23:0] _T_82639;
  wire [23:0] _GEN_7402;
  wire [23:0] _T_82643;
  wire [31:0] _GEN_7403;
  wire [31:0] _T_82679;
  wire [31:0] _GEN_7404;
  wire [31:0] _T_82683;
  wire [15:0] _GEN_7405;
  wire [15:0] _T_82759;
  wire [15:0] _GEN_7406;
  wire [15:0] _T_82763;
  wire [23:0] _GEN_7407;
  wire [23:0] _T_82799;
  wire [23:0] _GEN_7408;
  wire [23:0] _T_82803;
  wire [31:0] _GEN_7409;
  wire [31:0] _T_82839;
  wire [31:0] _GEN_7410;
  wire [31:0] _T_82843;
  wire  _T_82844;
  wire  _T_82845;
  wire  _T_82846;
  wire  _T_82847;
  wire  _T_82848;
  wire  _T_82849;
  wire  _T_82850;
  wire  _T_82851;
  wire  _T_82852;
  wire [1:0] _T_82854;
  wire [1:0] _T_82855;
  wire [3:0] _T_82856;
  wire [1:0] _T_82857;
  wire [1:0] _T_82858;
  wire [2:0] _T_82859;
  wire [4:0] _T_82860;
  wire [8:0] _T_82861;
  wire [511:0] _T_82881;
  wire  _T_82946;
  wire  _T_82947;
  wire  _T_82948;
  wire  _T_82949;
  wire  _T_83090;
  wire  _T_83091;
  wire  _T_83092;
  wire  _T_83093;
  wire  _T_83094;
  wire  _T_83095;
  wire  _T_83096;
  wire  _T_83097;
  wire  _T_83098;
  wire  _T_83099;
  wire  _T_83100;
  wire  _T_83101;
  wire  _T_83102;
  wire  _T_83103;
  wire  _T_83104;
  wire  _T_83105;
  wire  _T_83106;
  wire  _T_83908;
  wire  _T_88525;
  wire  _T_88526;
  wire  _T_89041;
  wire  _T_89049;
  wire  _T_89057;
  wire  _T_89065;
  wire  _T_90193;
  wire  _T_90201;
  wire  _T_90209;
  wire  _T_90217;
  wire  _T_90225;
  wire  _T_90233;
  wire  _T_90241;
  wire  _T_90249;
  wire  _T_90257;
  wire  _T_90265;
  wire  _T_90273;
  wire  _T_90281;
  wire  _T_90289;
  wire  _T_90297;
  wire  _T_90305;
  wire  _T_90313;
  wire  _T_90321;
  wire  _T_98274;
  wire  _T_98282;
  wire  _T_98290;
  wire  _T_98298;
  wire  _T_99426;
  wire  _T_99434;
  wire  _T_99442;
  wire  _T_99450;
  wire  _T_99458;
  wire  _T_99466;
  wire  _T_99474;
  wire  _T_99482;
  wire  _T_99490;
  wire  _T_99498;
  wire  _T_99506;
  wire  _T_99514;
  wire  _T_99522;
  wire  _T_99530;
  wire  _T_99538;
  wire  _T_99546;
  wire  _T_99554;
  wire [31:0] _T_102902_64;
  wire [31:0] _T_102902_65;
  wire [31:0] _T_102902_66;
  wire [31:0] _T_102902_67;
  wire  _GEN_4555;
  wire  _GEN_4556;
  wire  _GEN_4557;
  wire  _GEN_4558;
  wire  _GEN_4559;
  wire  _GEN_4560;
  wire  _GEN_4561;
  wire  _GEN_4562;
  wire  _GEN_4563;
  wire  _GEN_4564;
  wire  _GEN_4565;
  wire  _GEN_4566;
  wire  _GEN_4567;
  wire  _GEN_4568;
  wire  _GEN_4569;
  wire  _GEN_4570;
  wire  _GEN_4571;
  wire  _GEN_4572;
  wire  _GEN_4573;
  wire  _GEN_4574;
  wire  _GEN_4575;
  wire  _GEN_4576;
  wire  _GEN_4577;
  wire  _GEN_4578;
  wire  _GEN_4579;
  wire  _GEN_4580;
  wire  _GEN_4581;
  wire  _GEN_4582;
  wire  _GEN_4583;
  wire  _GEN_4584;
  wire  _GEN_4585;
  wire  _GEN_4586;
  wire  _GEN_4587;
  wire  _GEN_4588;
  wire  _GEN_4589;
  wire  _GEN_4590;
  wire  _GEN_4591;
  wire  _GEN_4592;
  wire  _GEN_4593;
  wire  _GEN_4594;
  wire  _GEN_4595;
  wire  _GEN_4596;
  wire  _GEN_4597;
  wire  _GEN_4598;
  wire  _GEN_4599;
  wire  _GEN_4600;
  wire  _GEN_4601;
  wire  _GEN_4602;
  wire  _GEN_4603;
  wire  _GEN_4604;
  wire  _GEN_4605;
  wire  _GEN_4606;
  wire  _GEN_4607;
  wire  _GEN_4608;
  wire  _GEN_4609;
  wire  _GEN_4610;
  wire  _GEN_4611;
  wire  _GEN_4612;
  wire  _GEN_4613;
  wire  _GEN_4614;
  wire  _GEN_4615;
  wire  _GEN_4616;
  wire  _GEN_4617;
  wire  _GEN_4618;
  wire  _GEN_4619;
  wire  _GEN_4620;
  wire  _GEN_4621;
  wire  _GEN_4622;
  wire  _GEN_4623;
  wire  _GEN_4624;
  wire  _GEN_4625;
  wire  _GEN_4626;
  wire  _GEN_4627;
  wire  _GEN_4628;
  wire  _GEN_4629;
  wire  _GEN_4630;
  wire  _GEN_4631;
  wire  _GEN_4632;
  wire  _GEN_4633;
  wire  _GEN_4634;
  wire  _GEN_4635;
  wire  _GEN_4636;
  wire  _GEN_4637;
  wire  _GEN_4638;
  wire  _GEN_4639;
  wire  _GEN_4640;
  wire  _GEN_4641;
  wire  _GEN_4642;
  wire  _GEN_4643;
  wire  _GEN_4644;
  wire  _GEN_4645;
  wire  _GEN_4646;
  wire  _GEN_4647;
  wire  _GEN_4648;
  wire  _GEN_4649;
  wire  _GEN_4650;
  wire  _GEN_4651;
  wire  _GEN_4652;
  wire  _GEN_4653;
  wire  _GEN_4654;
  wire  _GEN_4655;
  wire  _GEN_4656;
  wire  _GEN_4657;
  wire  _GEN_4658;
  wire  _GEN_4659;
  wire  _GEN_4660;
  wire  _GEN_4661;
  wire  _GEN_4662;
  wire  _GEN_4663;
  wire  _GEN_4664;
  wire  _GEN_4665;
  wire  _GEN_4666;
  wire  _GEN_4667;
  wire  _GEN_4668;
  wire  _GEN_4669;
  wire  _GEN_4670;
  wire  _GEN_4671;
  wire  _GEN_4672;
  wire  _GEN_4673;
  wire  _GEN_4674;
  wire  _GEN_4675;
  wire  _GEN_4676;
  wire  _GEN_4677;
  wire  _GEN_4678;
  wire  _GEN_4679;
  wire  _GEN_4680;
  wire  _GEN_4681;
  wire  _GEN_4682;
  wire  _GEN_4683;
  wire  _GEN_4684;
  wire  _GEN_4685;
  wire  _GEN_4686;
  wire  _GEN_4687;
  wire  _GEN_4688;
  wire  _GEN_4689;
  wire  _GEN_4690;
  wire  _GEN_4691;
  wire  _GEN_4692;
  wire  _GEN_4693;
  wire  _GEN_4694;
  wire  _GEN_4695;
  wire  _GEN_4696;
  wire  _GEN_4697;
  wire  _GEN_4698;
  wire  _GEN_4699;
  wire  _GEN_4700;
  wire  _GEN_4701;
  wire  _GEN_4702;
  wire  _GEN_4703;
  wire  _GEN_4704;
  wire  _GEN_4705;
  wire  _GEN_4706;
  wire  _GEN_4707;
  wire  _GEN_4708;
  wire  _GEN_4709;
  wire  _GEN_4710;
  wire  _GEN_4711;
  wire  _GEN_4712;
  wire  _GEN_4713;
  wire  _GEN_4714;
  wire  _GEN_4715;
  wire  _GEN_4716;
  wire  _GEN_4717;
  wire  _GEN_4718;
  wire  _GEN_4719;
  wire  _GEN_4720;
  wire  _GEN_4721;
  wire  _GEN_4722;
  wire  _GEN_4723;
  wire  _GEN_4724;
  wire  _GEN_4725;
  wire  _GEN_4726;
  wire  _GEN_4727;
  wire  _GEN_4728;
  wire  _GEN_4729;
  wire  _GEN_4730;
  wire  _GEN_4731;
  wire  _GEN_4732;
  wire  _GEN_4733;
  wire  _GEN_4734;
  wire  _GEN_4735;
  wire  _GEN_4736;
  wire  _GEN_4737;
  wire  _GEN_4738;
  wire  _GEN_4739;
  wire  _GEN_4740;
  wire  _GEN_4741;
  wire  _GEN_4742;
  wire  _GEN_4743;
  wire  _GEN_4744;
  wire  _GEN_4745;
  wire  _GEN_4746;
  wire  _GEN_4747;
  wire  _GEN_4748;
  wire  _GEN_4749;
  wire  _GEN_4750;
  wire  _GEN_4751;
  wire  _GEN_4752;
  wire  _GEN_4753;
  wire  _GEN_4754;
  wire  _GEN_4755;
  wire  _GEN_4756;
  wire  _GEN_4757;
  wire  _GEN_4758;
  wire  _GEN_4759;
  wire  _GEN_4760;
  wire  _GEN_4761;
  wire  _GEN_4762;
  wire  _GEN_4763;
  wire  _GEN_4764;
  wire  _GEN_4765;
  wire  _GEN_4766;
  wire  _GEN_4767;
  wire  _GEN_4768;
  wire  _GEN_4769;
  wire  _GEN_4770;
  wire  _GEN_4771;
  wire  _GEN_4772;
  wire  _GEN_4773;
  wire  _GEN_4774;
  wire  _GEN_4775;
  wire  _GEN_4776;
  wire  _GEN_4777;
  wire  _GEN_4778;
  wire  _GEN_4779;
  wire  _GEN_4780;
  wire  _GEN_4781;
  wire  _GEN_4782;
  wire  _GEN_4783;
  wire  _GEN_4784;
  wire  _GEN_4785;
  wire  _GEN_4786;
  wire  _GEN_4787;
  wire  _GEN_4788;
  wire  _GEN_4789;
  wire  _GEN_4790;
  wire  _GEN_4791;
  wire  _GEN_4792;
  wire  _GEN_4793;
  wire  _GEN_4794;
  wire  _GEN_4795;
  wire  _GEN_4796;
  wire  _GEN_4797;
  wire  _GEN_4798;
  wire  _GEN_4799;
  wire  _GEN_4800;
  wire  _GEN_4801;
  wire  _GEN_4802;
  wire  _GEN_4803;
  wire  _GEN_4804;
  wire  _GEN_4805;
  wire  _GEN_4806;
  wire  _GEN_4807;
  wire  _GEN_4808;
  wire  _GEN_4809;
  wire  _GEN_4810;
  wire  _GEN_4811;
  wire  _GEN_4812;
  wire  _GEN_4813;
  wire  _GEN_4814;
  wire  _GEN_4815;
  wire  _GEN_4816;
  wire  _GEN_4817;
  wire  _GEN_4818;
  wire  _GEN_4819;
  wire  _GEN_4820;
  wire  _GEN_4821;
  wire  _GEN_4822;
  wire  _GEN_4823;
  wire  _GEN_4824;
  wire  _GEN_4825;
  wire  _GEN_4826;
  wire  _GEN_4827;
  wire  _GEN_4828;
  wire  _GEN_4829;
  wire  _GEN_4830;
  wire  _GEN_4831;
  wire  _GEN_4832;
  wire  _GEN_4833;
  wire  _GEN_4834;
  wire  _GEN_4835;
  wire  _GEN_4836;
  wire  _GEN_4837;
  wire  _GEN_4838;
  wire  _GEN_4839;
  wire  _GEN_4840;
  wire  _GEN_4841;
  wire  _GEN_4842;
  wire  _GEN_4843;
  wire  _GEN_4844;
  wire  _GEN_4845;
  wire  _GEN_4846;
  wire  _GEN_4847;
  wire  _GEN_4848;
  wire  _GEN_4849;
  wire  _GEN_4850;
  wire  _GEN_4851;
  wire  _GEN_4852;
  wire  _GEN_4853;
  wire  _GEN_4854;
  wire  _GEN_4855;
  wire  _GEN_4856;
  wire  _GEN_4857;
  wire  _GEN_4858;
  wire  _GEN_4859;
  wire  _GEN_4860;
  wire  _GEN_4861;
  wire  _GEN_4862;
  wire  _GEN_4863;
  wire  _GEN_4864;
  wire  _GEN_4865;
  wire  _GEN_4866;
  wire  _GEN_4867;
  wire  _GEN_4868;
  wire  _GEN_4869;
  wire  _GEN_4870;
  wire  _GEN_4871;
  wire  _GEN_4872;
  wire  _GEN_4873;
  wire  _GEN_4874;
  wire  _GEN_4875;
  wire  _GEN_4876;
  wire  _GEN_4877;
  wire  _GEN_4878;
  wire  _GEN_4879;
  wire  _GEN_4880;
  wire  _GEN_4881;
  wire  _GEN_4882;
  wire  _GEN_4883;
  wire  _GEN_4884;
  wire  _GEN_4885;
  wire  _GEN_4886;
  wire  _GEN_4887;
  wire  _GEN_4888;
  wire  _GEN_4889;
  wire  _GEN_4890;
  wire  _GEN_4891;
  wire  _GEN_4892;
  wire  _GEN_4893;
  wire  _GEN_4894;
  wire  _GEN_4895;
  wire  _GEN_4896;
  wire  _GEN_4897;
  wire  _GEN_4898;
  wire  _GEN_4899;
  wire  _GEN_4900;
  wire  _GEN_4901;
  wire  _GEN_4902;
  wire  _GEN_4903;
  wire  _GEN_4904;
  wire  _GEN_4905;
  wire  _GEN_4906;
  wire  _GEN_4907;
  wire  _GEN_4908;
  wire  _GEN_4909;
  wire  _GEN_4910;
  wire  _GEN_4911;
  wire  _GEN_4912;
  wire  _GEN_4913;
  wire  _GEN_4914;
  wire  _GEN_4915;
  wire  _GEN_4916;
  wire  _GEN_4917;
  wire  _GEN_4918;
  wire  _GEN_4919;
  wire  _GEN_4920;
  wire  _GEN_4921;
  wire  _GEN_4922;
  wire  _GEN_4923;
  wire  _GEN_4924;
  wire  _GEN_4925;
  wire  _GEN_4926;
  wire  _GEN_4927;
  wire  _GEN_4928;
  wire  _GEN_4929;
  wire  _GEN_4930;
  wire  _GEN_4931;
  wire  _GEN_4932;
  wire  _GEN_4933;
  wire  _GEN_4934;
  wire  _GEN_4935;
  wire  _GEN_4936;
  wire  _GEN_4937;
  wire  _GEN_4938;
  wire  _GEN_4939;
  wire  _GEN_4940;
  wire  _GEN_4941;
  wire  _GEN_4942;
  wire  _GEN_4943;
  wire  _GEN_4944;
  wire  _GEN_4945;
  wire  _GEN_4946;
  wire  _GEN_4947;
  wire  _GEN_4948;
  wire  _GEN_4949;
  wire  _GEN_4950;
  wire  _GEN_4951;
  wire  _GEN_4952;
  wire  _GEN_4953;
  wire  _GEN_4954;
  wire  _GEN_4955;
  wire  _GEN_4956;
  wire  _GEN_4957;
  wire  _GEN_4958;
  wire  _GEN_4959;
  wire  _GEN_4960;
  wire  _GEN_4961;
  wire  _GEN_4962;
  wire  _GEN_4963;
  wire  _GEN_4964;
  wire  _GEN_4965;
  wire  _GEN_4966;
  wire  _GEN_4967;
  wire  _GEN_4968;
  wire  _GEN_4969;
  wire  _GEN_4970;
  wire  _GEN_4971;
  wire  _GEN_4972;
  wire  _GEN_4973;
  wire  _GEN_4974;
  wire  _GEN_4975;
  wire  _GEN_4976;
  wire  _GEN_4977;
  wire  _GEN_4978;
  wire  _GEN_4979;
  wire  _GEN_4980;
  wire  _GEN_4981;
  wire  _GEN_4982;
  wire  _GEN_4983;
  wire  _GEN_4984;
  wire  _GEN_4985;
  wire  _GEN_4986;
  wire  _GEN_4987;
  wire  _GEN_4988;
  wire  _GEN_4989;
  wire  _GEN_4990;
  wire  _GEN_4991;
  wire  _GEN_4992;
  wire  _GEN_4993;
  wire  _GEN_4994;
  wire  _GEN_4995;
  wire  _GEN_4996;
  wire  _GEN_4997;
  wire  _GEN_4998;
  wire  _GEN_4999;
  wire  _GEN_5000;
  wire  _GEN_5001;
  wire  _GEN_5002;
  wire  _GEN_5003;
  wire  _GEN_5004;
  wire  _GEN_5005;
  wire  _GEN_5006;
  wire  _GEN_5007;
  wire  _GEN_5008;
  wire  _GEN_5009;
  wire  _GEN_5010;
  wire  _GEN_5011;
  wire  _GEN_5012;
  wire  _GEN_5013;
  wire  _GEN_5014;
  wire  _GEN_5015;
  wire  _GEN_5016;
  wire  _GEN_5017;
  wire  _GEN_5018;
  wire  _GEN_5019;
  wire  _GEN_5020;
  wire  _GEN_5021;
  wire  _GEN_5022;
  wire  _GEN_5023;
  wire  _GEN_5024;
  wire  _GEN_5025;
  wire  _GEN_5026;
  wire  _GEN_5027;
  wire  _GEN_5028;
  wire  _GEN_5029;
  wire  _GEN_5030;
  wire  _GEN_5031;
  wire  _GEN_5032;
  wire  _GEN_5033;
  wire  _GEN_5034;
  wire  _GEN_5035;
  wire  _GEN_5036;
  wire  _GEN_5037;
  wire  _GEN_5038;
  wire  _GEN_5039;
  wire  _GEN_5040;
  wire  _GEN_5041;
  wire  _GEN_5042;
  wire  _GEN_5043;
  wire  _GEN_5044;
  wire  _GEN_5045;
  wire  _GEN_5046;
  wire  _GEN_5047;
  wire  _GEN_5048;
  wire  _GEN_5049;
  wire  _GEN_5050;
  wire  _GEN_5051;
  wire  _GEN_5052;
  wire  _GEN_5053;
  wire  _GEN_5054;
  wire  _GEN_5055;
  wire  _GEN_5056;
  wire  _GEN_5057;
  wire  _GEN_5058;
  wire  _GEN_5059;
  wire  _GEN_5060;
  wire  _GEN_5061;
  wire  _GEN_5062;
  wire  _GEN_5063;
  wire  _GEN_5064;
  wire  _GEN_5065;
  wire [31:0] _GEN_5066;
  wire [31:0] _GEN_5067;
  wire [31:0] _GEN_5068;
  wire [31:0] _GEN_5069;
  wire [31:0] _GEN_5070;
  wire [31:0] _GEN_5071;
  wire [31:0] _GEN_5072;
  wire [31:0] _GEN_5073;
  wire [31:0] _GEN_5074;
  wire [31:0] _GEN_5075;
  wire [31:0] _GEN_5076;
  wire [31:0] _GEN_5077;
  wire [31:0] _GEN_5078;
  wire [31:0] _GEN_5079;
  wire [31:0] _GEN_5080;
  wire [31:0] _GEN_5081;
  wire [31:0] _GEN_5082;
  wire [31:0] _GEN_5083;
  wire [31:0] _GEN_5084;
  wire [31:0] _GEN_5085;
  wire [31:0] _GEN_5086;
  wire [31:0] _GEN_5087;
  wire [31:0] _GEN_5088;
  wire [31:0] _GEN_5089;
  wire [31:0] _GEN_5090;
  wire [31:0] _GEN_5091;
  wire [31:0] _GEN_5092;
  wire [31:0] _GEN_5093;
  wire [31:0] _GEN_5094;
  wire [31:0] _GEN_5095;
  wire [31:0] _GEN_5096;
  wire [31:0] _GEN_5097;
  wire [31:0] _GEN_5098;
  wire [31:0] _GEN_5099;
  wire [31:0] _GEN_5100;
  wire [31:0] _GEN_5101;
  wire [31:0] _GEN_5102;
  wire [31:0] _GEN_5103;
  wire [31:0] _GEN_5104;
  wire [31:0] _GEN_5105;
  wire [31:0] _GEN_5106;
  wire [31:0] _GEN_5107;
  wire [31:0] _GEN_5108;
  wire [31:0] _GEN_5109;
  wire [31:0] _GEN_5110;
  wire [31:0] _GEN_5111;
  wire [31:0] _GEN_5112;
  wire [31:0] _GEN_5113;
  wire [31:0] _GEN_5114;
  wire [31:0] _GEN_5115;
  wire [31:0] _GEN_5116;
  wire [31:0] _GEN_5117;
  wire [31:0] _GEN_5118;
  wire [31:0] _GEN_5119;
  wire [31:0] _GEN_5120;
  wire [31:0] _GEN_5121;
  wire [31:0] _GEN_5122;
  wire [31:0] _GEN_5123;
  wire [31:0] _GEN_5124;
  wire [31:0] _GEN_5125;
  wire [31:0] _GEN_5126;
  wire [31:0] _GEN_5127;
  wire [31:0] _GEN_5128;
  wire [31:0] _GEN_5129;
  wire [31:0] _GEN_5130;
  wire [31:0] _GEN_5131;
  wire [31:0] _GEN_5132;
  wire [31:0] _GEN_5133;
  wire [31:0] _GEN_5134;
  wire [31:0] _GEN_5135;
  wire [31:0] _GEN_5136;
  wire [31:0] _GEN_5137;
  wire [31:0] _GEN_5138;
  wire [31:0] _GEN_5139;
  wire [31:0] _GEN_5140;
  wire [31:0] _GEN_5141;
  wire [31:0] _GEN_5142;
  wire [31:0] _GEN_5143;
  wire [31:0] _GEN_5144;
  wire [31:0] _GEN_5145;
  wire [31:0] _GEN_5146;
  wire [31:0] _GEN_5147;
  wire [31:0] _GEN_5148;
  wire [31:0] _GEN_5149;
  wire [31:0] _GEN_5150;
  wire [31:0] _GEN_5151;
  wire [31:0] _GEN_5152;
  wire [31:0] _GEN_5153;
  wire [31:0] _GEN_5154;
  wire [31:0] _GEN_5155;
  wire [31:0] _GEN_5156;
  wire [31:0] _GEN_5157;
  wire [31:0] _GEN_5158;
  wire [31:0] _GEN_5159;
  wire [31:0] _GEN_5160;
  wire [31:0] _GEN_5161;
  wire [31:0] _GEN_5162;
  wire [31:0] _GEN_5163;
  wire [31:0] _GEN_5164;
  wire [31:0] _GEN_5165;
  wire [31:0] _GEN_5166;
  wire [31:0] _GEN_5167;
  wire [31:0] _GEN_5168;
  wire [31:0] _GEN_5169;
  wire [31:0] _GEN_5170;
  wire [31:0] _GEN_5171;
  wire [31:0] _GEN_5172;
  wire [31:0] _GEN_5173;
  wire [31:0] _GEN_5174;
  wire [31:0] _GEN_5175;
  wire [31:0] _GEN_5176;
  wire [31:0] _GEN_5177;
  wire [31:0] _GEN_5178;
  wire [31:0] _GEN_5179;
  wire [31:0] _GEN_5180;
  wire [31:0] _GEN_5181;
  wire [31:0] _GEN_5182;
  wire [31:0] _GEN_5183;
  wire [31:0] _GEN_5184;
  wire [31:0] _GEN_5185;
  wire [31:0] _GEN_5186;
  wire [31:0] _GEN_5187;
  wire [31:0] _GEN_5188;
  wire [31:0] _GEN_5189;
  wire [31:0] _GEN_5190;
  wire [31:0] _GEN_5191;
  wire [31:0] _GEN_5192;
  wire [31:0] _GEN_5193;
  wire [31:0] _GEN_5194;
  wire [31:0] _GEN_5195;
  wire [31:0] _GEN_5196;
  wire [31:0] _GEN_5197;
  wire [31:0] _GEN_5198;
  wire [31:0] _GEN_5199;
  wire [31:0] _GEN_5200;
  wire [31:0] _GEN_5201;
  wire [31:0] _GEN_5202;
  wire [31:0] _GEN_5203;
  wire [31:0] _GEN_5204;
  wire [31:0] _GEN_5205;
  wire [31:0] _GEN_5206;
  wire [31:0] _GEN_5207;
  wire [31:0] _GEN_5208;
  wire [31:0] _GEN_5209;
  wire [31:0] _GEN_5210;
  wire [31:0] _GEN_5211;
  wire [31:0] _GEN_5212;
  wire [31:0] _GEN_5213;
  wire [31:0] _GEN_5214;
  wire [31:0] _GEN_5215;
  wire [31:0] _GEN_5216;
  wire [31:0] _GEN_5217;
  wire [31:0] _GEN_5218;
  wire [31:0] _GEN_5219;
  wire [31:0] _GEN_5220;
  wire [31:0] _GEN_5221;
  wire [31:0] _GEN_5222;
  wire [31:0] _GEN_5223;
  wire [31:0] _GEN_5224;
  wire [31:0] _GEN_5225;
  wire [31:0] _GEN_5226;
  wire [31:0] _GEN_5227;
  wire [31:0] _GEN_5228;
  wire [31:0] _GEN_5229;
  wire [31:0] _GEN_5230;
  wire [31:0] _GEN_5231;
  wire [31:0] _GEN_5232;
  wire [31:0] _GEN_5233;
  wire [31:0] _GEN_5234;
  wire [31:0] _GEN_5235;
  wire [31:0] _GEN_5236;
  wire [31:0] _GEN_5237;
  wire [31:0] _GEN_5238;
  wire [31:0] _GEN_5239;
  wire [31:0] _GEN_5240;
  wire [31:0] _GEN_5241;
  wire [31:0] _GEN_5242;
  wire [31:0] _GEN_5243;
  wire [31:0] _GEN_5244;
  wire [31:0] _GEN_5245;
  wire [31:0] _GEN_5246;
  wire [31:0] _GEN_5247;
  wire [31:0] _GEN_5248;
  wire [31:0] _GEN_5249;
  wire [31:0] _GEN_5250;
  wire [31:0] _GEN_5251;
  wire [31:0] _GEN_5252;
  wire [31:0] _GEN_5253;
  wire [31:0] _GEN_5254;
  wire [31:0] _GEN_5255;
  wire [31:0] _GEN_5256;
  wire [31:0] _GEN_5257;
  wire [31:0] _GEN_5258;
  wire [31:0] _GEN_5259;
  wire [31:0] _GEN_5260;
  wire [31:0] _GEN_5261;
  wire [31:0] _GEN_5262;
  wire [31:0] _GEN_5263;
  wire [31:0] _GEN_5264;
  wire [31:0] _GEN_5265;
  wire [31:0] _GEN_5266;
  wire [31:0] _GEN_5267;
  wire [31:0] _GEN_5268;
  wire [31:0] _GEN_5269;
  wire [31:0] _GEN_5270;
  wire [31:0] _GEN_5271;
  wire [31:0] _GEN_5272;
  wire [31:0] _GEN_5273;
  wire [31:0] _GEN_5274;
  wire [31:0] _GEN_5275;
  wire [31:0] _GEN_5276;
  wire [31:0] _GEN_5277;
  wire [31:0] _GEN_5278;
  wire [31:0] _GEN_5279;
  wire [31:0] _GEN_5280;
  wire [31:0] _GEN_5281;
  wire [31:0] _GEN_5282;
  wire [31:0] _GEN_5283;
  wire [31:0] _GEN_5284;
  wire [31:0] _GEN_5285;
  wire [31:0] _GEN_5286;
  wire [31:0] _GEN_5287;
  wire [31:0] _GEN_5288;
  wire [31:0] _GEN_5289;
  wire [31:0] _GEN_5290;
  wire [31:0] _GEN_5291;
  wire [31:0] _GEN_5292;
  wire [31:0] _GEN_5293;
  wire [31:0] _GEN_5294;
  wire [31:0] _GEN_5295;
  wire [31:0] _GEN_5296;
  wire [31:0] _GEN_5297;
  wire [31:0] _GEN_5298;
  wire [31:0] _GEN_5299;
  wire [31:0] _GEN_5300;
  wire [31:0] _GEN_5301;
  wire [31:0] _GEN_5302;
  wire [31:0] _GEN_5303;
  wire [31:0] _GEN_5304;
  wire [31:0] _GEN_5305;
  wire [31:0] _GEN_5306;
  wire [31:0] _GEN_5307;
  wire [31:0] _GEN_5308;
  wire [31:0] _GEN_5309;
  wire [31:0] _GEN_5310;
  wire [31:0] _GEN_5311;
  wire [31:0] _GEN_5312;
  wire [31:0] _GEN_5313;
  wire [31:0] _GEN_5314;
  wire [31:0] _GEN_5315;
  wire [31:0] _GEN_5316;
  wire [31:0] _GEN_5317;
  wire [31:0] _GEN_5318;
  wire [31:0] _GEN_5319;
  wire [31:0] _GEN_5320;
  wire [31:0] _GEN_5321;
  wire [31:0] _GEN_5322;
  wire [31:0] _GEN_5323;
  wire [31:0] _GEN_5324;
  wire [31:0] _GEN_5325;
  wire [31:0] _GEN_5326;
  wire [31:0] _GEN_5327;
  wire [31:0] _GEN_5328;
  wire [31:0] _GEN_5329;
  wire [31:0] _GEN_5330;
  wire [31:0] _GEN_5331;
  wire [31:0] _GEN_5332;
  wire [31:0] _GEN_5333;
  wire [31:0] _GEN_5334;
  wire [31:0] _GEN_5335;
  wire [31:0] _GEN_5336;
  wire [31:0] _GEN_5337;
  wire [31:0] _GEN_5338;
  wire [31:0] _GEN_5339;
  wire [31:0] _GEN_5340;
  wire [31:0] _GEN_5341;
  wire [31:0] _GEN_5342;
  wire [31:0] _GEN_5343;
  wire [31:0] _GEN_5344;
  wire [31:0] _GEN_5345;
  wire [31:0] _GEN_5346;
  wire [31:0] _GEN_5347;
  wire [31:0] _GEN_5348;
  wire [31:0] _GEN_5349;
  wire [31:0] _GEN_5350;
  wire [31:0] _GEN_5351;
  wire [31:0] _GEN_5352;
  wire [31:0] _GEN_5353;
  wire [31:0] _GEN_5354;
  wire [31:0] _GEN_5355;
  wire [31:0] _GEN_5356;
  wire [31:0] _GEN_5357;
  wire [31:0] _GEN_5358;
  wire [31:0] _GEN_5359;
  wire [31:0] _GEN_5360;
  wire [31:0] _GEN_5361;
  wire [31:0] _GEN_5362;
  wire [31:0] _GEN_5363;
  wire [31:0] _GEN_5364;
  wire [31:0] _GEN_5365;
  wire [31:0] _GEN_5366;
  wire [31:0] _GEN_5367;
  wire [31:0] _GEN_5368;
  wire [31:0] _GEN_5369;
  wire [31:0] _GEN_5370;
  wire [31:0] _GEN_5371;
  wire [31:0] _GEN_5372;
  wire [31:0] _GEN_5373;
  wire [31:0] _GEN_5374;
  wire [31:0] _GEN_5375;
  wire [31:0] _GEN_5376;
  wire [31:0] _GEN_5377;
  wire [31:0] _GEN_5378;
  wire [31:0] _GEN_5379;
  wire [31:0] _GEN_5380;
  wire [31:0] _GEN_5381;
  wire [31:0] _GEN_5382;
  wire [31:0] _GEN_5383;
  wire [31:0] _GEN_5384;
  wire [31:0] _GEN_5385;
  wire [31:0] _GEN_5386;
  wire [31:0] _GEN_5387;
  wire [31:0] _GEN_5388;
  wire [31:0] _GEN_5389;
  wire [31:0] _GEN_5390;
  wire [31:0] _GEN_5391;
  wire [31:0] _GEN_5392;
  wire [31:0] _GEN_5393;
  wire [31:0] _GEN_5394;
  wire [31:0] _GEN_5395;
  wire [31:0] _GEN_5396;
  wire [31:0] _GEN_5397;
  wire [31:0] _GEN_5398;
  wire [31:0] _GEN_5399;
  wire [31:0] _GEN_5400;
  wire [31:0] _GEN_5401;
  wire [31:0] _GEN_5402;
  wire [31:0] _GEN_5403;
  wire [31:0] _GEN_5404;
  wire [31:0] _GEN_5405;
  wire [31:0] _GEN_5406;
  wire [31:0] _GEN_5407;
  wire [31:0] _GEN_5408;
  wire [31:0] _GEN_5409;
  wire [31:0] _GEN_5410;
  wire [31:0] _GEN_5411;
  wire [31:0] _GEN_5412;
  wire [31:0] _GEN_5413;
  wire [31:0] _GEN_5414;
  wire [31:0] _GEN_5415;
  wire [31:0] _GEN_5416;
  wire [31:0] _GEN_5417;
  wire [31:0] _GEN_5418;
  wire [31:0] _GEN_5419;
  wire [31:0] _GEN_5420;
  wire [31:0] _GEN_5421;
  wire [31:0] _GEN_5422;
  wire [31:0] _GEN_5423;
  wire [31:0] _GEN_5424;
  wire [31:0] _GEN_5425;
  wire [31:0] _GEN_5426;
  wire [31:0] _GEN_5427;
  wire [31:0] _GEN_5428;
  wire [31:0] _GEN_5429;
  wire [31:0] _GEN_5430;
  wire [31:0] _GEN_5431;
  wire [31:0] _GEN_5432;
  wire [31:0] _GEN_5433;
  wire [31:0] _GEN_5434;
  wire [31:0] _GEN_5435;
  wire [31:0] _GEN_5436;
  wire [31:0] _GEN_5437;
  wire [31:0] _GEN_5438;
  wire [31:0] _GEN_5439;
  wire [31:0] _GEN_5440;
  wire [31:0] _GEN_5441;
  wire [31:0] _GEN_5442;
  wire [31:0] _GEN_5443;
  wire [31:0] _GEN_5444;
  wire [31:0] _GEN_5445;
  wire [31:0] _GEN_5446;
  wire [31:0] _GEN_5447;
  wire [31:0] _GEN_5448;
  wire [31:0] _GEN_5449;
  wire [31:0] _GEN_5450;
  wire [31:0] _GEN_5451;
  wire [31:0] _GEN_5452;
  wire [31:0] _GEN_5453;
  wire [31:0] _GEN_5454;
  wire [31:0] _GEN_5455;
  wire [31:0] _GEN_5456;
  wire [31:0] _GEN_5457;
  wire [31:0] _GEN_5458;
  wire [31:0] _GEN_5459;
  wire [31:0] _GEN_5460;
  wire [31:0] _GEN_5461;
  wire [31:0] _GEN_5462;
  wire [31:0] _GEN_5463;
  wire [31:0] _GEN_5464;
  wire [31:0] _GEN_5465;
  wire [31:0] _GEN_5466;
  wire [31:0] _GEN_5467;
  wire [31:0] _GEN_5468;
  wire [31:0] _GEN_5469;
  wire [31:0] _GEN_5470;
  wire [31:0] _GEN_5471;
  wire [31:0] _GEN_5472;
  wire [31:0] _GEN_5473;
  wire [31:0] _GEN_5474;
  wire [31:0] _GEN_5475;
  wire [31:0] _GEN_5476;
  wire [31:0] _GEN_5477;
  wire [31:0] _GEN_5478;
  wire [31:0] _GEN_5479;
  wire [31:0] _GEN_5480;
  wire [31:0] _GEN_5481;
  wire [31:0] _GEN_5482;
  wire [31:0] _GEN_5483;
  wire [31:0] _GEN_5484;
  wire [31:0] _GEN_5485;
  wire [31:0] _GEN_5486;
  wire [31:0] _GEN_5487;
  wire [31:0] _GEN_5488;
  wire [31:0] _GEN_5489;
  wire [31:0] _GEN_5490;
  wire [31:0] _GEN_5491;
  wire [31:0] _GEN_5492;
  wire [31:0] _GEN_5493;
  wire [31:0] _GEN_5494;
  wire [31:0] _GEN_5495;
  wire [31:0] _GEN_5496;
  wire [31:0] _GEN_5497;
  wire [31:0] _GEN_5498;
  wire [31:0] _GEN_5499;
  wire [31:0] _GEN_5500;
  wire [31:0] _GEN_5501;
  wire [31:0] _GEN_5502;
  wire [31:0] _GEN_5503;
  wire [31:0] _GEN_5504;
  wire [31:0] _GEN_5505;
  wire [31:0] _GEN_5506;
  wire [31:0] _GEN_5507;
  wire [31:0] _GEN_5508;
  wire [31:0] _GEN_5509;
  wire [31:0] _GEN_5510;
  wire [31:0] _GEN_5511;
  wire [31:0] _GEN_5512;
  wire [31:0] _GEN_5513;
  wire [31:0] _GEN_5514;
  wire [31:0] _GEN_5515;
  wire [31:0] _GEN_5516;
  wire [31:0] _GEN_5517;
  wire [31:0] _GEN_5518;
  wire [31:0] _GEN_5519;
  wire [31:0] _GEN_5520;
  wire [31:0] _GEN_5521;
  wire [31:0] _GEN_5522;
  wire [31:0] _GEN_5523;
  wire [31:0] _GEN_5524;
  wire [31:0] _GEN_5525;
  wire [31:0] _GEN_5526;
  wire [31:0] _GEN_5527;
  wire [31:0] _GEN_5528;
  wire [31:0] _GEN_5529;
  wire [31:0] _GEN_5530;
  wire [31:0] _GEN_5531;
  wire [31:0] _GEN_5532;
  wire [31:0] _GEN_5533;
  wire [31:0] _GEN_5534;
  wire [31:0] _GEN_5535;
  wire [31:0] _GEN_5536;
  wire [31:0] _GEN_5537;
  wire [31:0] _GEN_5538;
  wire [31:0] _GEN_5539;
  wire [31:0] _GEN_5540;
  wire [31:0] _GEN_5541;
  wire [31:0] _GEN_5542;
  wire [31:0] _GEN_5543;
  wire [31:0] _GEN_5544;
  wire [31:0] _GEN_5545;
  wire [31:0] _GEN_5546;
  wire [31:0] _GEN_5547;
  wire [31:0] _GEN_5548;
  wire [31:0] _GEN_5549;
  wire [31:0] _GEN_5550;
  wire [31:0] _GEN_5551;
  wire [31:0] _GEN_5552;
  wire [31:0] _GEN_5553;
  wire [31:0] _GEN_5554;
  wire [31:0] _GEN_5555;
  wire [31:0] _GEN_5556;
  wire [31:0] _GEN_5557;
  wire [31:0] _GEN_5558;
  wire [31:0] _GEN_5559;
  wire [31:0] _GEN_5560;
  wire [31:0] _GEN_5561;
  wire [31:0] _GEN_5562;
  wire [31:0] _GEN_5563;
  wire [31:0] _GEN_5564;
  wire [31:0] _GEN_5565;
  wire [31:0] _GEN_5566;
  wire [31:0] _GEN_5567;
  wire [31:0] _GEN_5568;
  wire [31:0] _GEN_5569;
  wire [31:0] _GEN_5570;
  wire [31:0] _GEN_5571;
  wire [31:0] _GEN_5572;
  wire [31:0] _GEN_5573;
  wire [31:0] _GEN_5574;
  wire [31:0] _GEN_5575;
  wire [31:0] _GEN_5576;
  wire [31:0] _T_103419;
  wire [9:0] _T_103420;
  wire [1:0] _T_103421;
  wire [7:0] _GEN_5577;
  wire [7:0] _GEN_5578;
  wire [7:0] _GEN_5579;
  wire [7:0] _GEN_5580;
  wire [7:0] _GEN_5581;
  wire [7:0] _GEN_5582;
  wire [7:0] _GEN_5583;
  wire [7:0] _GEN_5584;
  wire [7:0] _GEN_5585;
  wire [7:0] _GEN_5586;
  wire [7:0] _GEN_5587;
  wire [7:0] _GEN_5588;
  wire [7:0] _GEN_5589;
  wire [7:0] _GEN_5590;
  wire [7:0] _GEN_5591;
  wire [7:0] _GEN_5592;
  wire [7:0] _GEN_5593;
  wire [7:0] _GEN_5594;
  wire [7:0] _GEN_5595;
  wire [7:0] _GEN_5596;
  wire [7:0] _GEN_5597;
  wire [7:0] _GEN_5598;
  wire [7:0] _GEN_5599;
  wire [7:0] _GEN_5600;
  wire [7:0] _GEN_5601;
  wire [7:0] _GEN_5602;
  wire [7:0] _GEN_5603;
  wire [7:0] _GEN_5604;
  wire [7:0] _GEN_5605;
  wire [7:0] _GEN_5606;
  wire [7:0] _GEN_5607;
  wire [7:0] _GEN_5608;
  wire [7:0] _GEN_5609;
  wire [7:0] _GEN_5610;
  wire [7:0] _GEN_5611;
  wire [7:0] _GEN_5612;
  wire [7:0] _GEN_5613;
  wire [7:0] _GEN_5614;
  wire [7:0] _GEN_5615;
  wire [7:0] _GEN_5616;
  wire [7:0] _GEN_5617;
  wire [7:0] _GEN_5618;
  wire [7:0] _GEN_5619;
  wire [7:0] _GEN_5620;
  wire [7:0] _GEN_5621;
  wire [7:0] _GEN_5622;
  wire [7:0] _GEN_5623;
  wire [7:0] _GEN_5624;
  wire [7:0] _GEN_5625;
  wire [7:0] _GEN_5626;
  wire [7:0] _GEN_5627;
  wire [7:0] _GEN_5628;
  wire [7:0] _GEN_5629;
  wire [7:0] _GEN_5630;
  wire [7:0] _GEN_5631;
  wire [7:0] _GEN_5632;
  wire [7:0] _GEN_5633;
  wire [7:0] _GEN_5634;
  wire [7:0] _GEN_5635;
  wire [7:0] _GEN_5636;
  wire [7:0] _GEN_5637;
  wire [7:0] _GEN_5638;
  wire [7:0] _GEN_5639;
  wire [7:0] _GEN_5640;
  wire [7:0] _GEN_5641;
  wire [7:0] _GEN_5642;
  wire [7:0] _GEN_5643;
  wire [7:0] _GEN_5644;
  reg [1:0] ctrlStateReg;
  reg [31:0] _RAND_86;
  wire  _T_103511;
  wire  _T_103513;
  wire  _T_103515;
  wire  _T_103517;
  wire  _T_103519;
  wire  _T_103521;
  wire  _T_103522;
  wire  _T_103523;
  wire  _T_103525;
  wire  _T_103526;
  wire  _T_103528;
  wire  _T_103529;
  wire  _T_103531;
  wire  _T_103532;
  wire  _T_103534;
  wire  _T_103535;
  wire  commandWrIsAccessRegister;
  wire  commandRegIsAccessRegister;
  wire  _T_103539;
  wire  commandWrIsUnsupported;
  wire  _T_103545;
  wire  _T_103547;
  wire  _T_103549;
  wire  _T_103550;
  wire  _T_103551;
  wire  _T_103553;
  wire  _GEN_5645;
  wire  _GEN_5646;
  wire  _GEN_5647;
  wire  _GEN_5648;
  wire  _T_103554;
  wire  _T_103556;
  wire  wrAccessRegisterCommand;
  wire  _T_103557;
  wire  regAccessRegisterCommand;
  wire  _T_103562;
  wire [1:0] _GEN_5649;
  wire  _T_103565;
  wire  _T_103566;
  wire  _T_103568;
  wire  _T_103572;
  wire  _T_103573;
  wire  _T_103574;
  wire  _GEN_5651;
  wire [1:0] _GEN_5652;
  wire  _GEN_5653;
  wire  _T_103577;
  wire  _T_103579;
  wire  _T_103580;
  wire  _GEN_5654;
  wire [1:0] _GEN_5655;
  wire  _T_103584;
  wire  _T_103585;
  wire [1:0] _GEN_5657;
  wire  _T_103591;
  wire  _T_103592;
  wire [1:0] _GEN_5658;
  wire  _GEN_5660;
  wire [1:0] _GEN_5661;
  wire  _GEN_5662;
  wire  _GEN_5663;
  wire  _T_103596;
  wire  _T_103600;
  wire  _T_103601;
  wire  _T_103602;
  wire  _T_103604;
  wire  _T_103605;
  wire  _T_103606;
  wire  _T_103607;
  wire [1:0] _GEN_5664;
  wire [1:0] _GEN_5665;
  wire [1:0] _GEN_5667;
  wire  _GEN_5668;
  wire [1:0] _GEN_5669;
  wire [1:0] _GEN_5670;
  wire  _GEN_7411;
  wire  _GEN_7413;
  assign io_hart_in_0_a_ready = io_hart_in_0_d_ready;
  assign io_hart_in_0_d_valid = io_hart_in_0_a_valid;
  assign io_hart_in_0_d_bits_opcode = {{2'd0}, _T_25899};
  assign io_hart_in_0_d_bits_param = 2'h0;
  assign io_hart_in_0_d_bits_size = _T_103421;
  assign io_hart_in_0_d_bits_source = _T_103420;
  assign io_hart_in_0_d_bits_sink = 1'h0;
  assign io_hart_in_0_d_bits_data = _T_103419;
  assign io_hart_in_0_d_bits_error = 1'h0;
  assign io_dmi_in_0_a_ready = io_dmi_in_0_d_ready;
  assign io_dmi_in_0_d_valid = io_dmi_in_0_a_valid;
  assign io_dmi_in_0_d_bits_opcode = {{2'd0}, _T_2874};
  assign io_dmi_in_0_d_bits_param = 2'h0;
  assign io_dmi_in_0_d_bits_size = _T_7942;
  assign io_dmi_in_0_d_bits_source = _T_7941;
  assign io_dmi_in_0_d_bits_sink = 1'h0;
  assign io_dmi_in_0_d_bits_data = _T_7940;
  assign io_dmi_in_0_d_bits_error = 1'h0;
  assign io_innerCtrl_ready = 1'h1;
  assign _T_1197 = io_innerCtrl_ready & io_innerCtrl_valid;
  assign _GEN_14 = _T_1197 ? io_innerCtrl_bits_hartsel : selectedHartReg;
  assign _T_1246 = selectedHartReg >= 10'h1;
  assign _T_1254 = _T_1246 == 1'h0;
  assign _T_1255 = _T_1254 & io_debugUnavail_0;
  assign _T_1265 = io_debugUnavail_0 == 1'h0;
  assign _T_1266 = _T_1254 & _T_1265;
  assign _T_1267 = _T_1266 & haltedBitRegs_0;
  assign _T_1276 = haltedBitRegs_0 == 1'h0;
  assign _T_1277 = _T_1266 & _T_1276;
  assign resumereq = _T_1197 & io_innerCtrl_bits_resumereq;
  assign _T_1285 = ~ resumeReqRegs_0;
  assign _T_1286 = ~ resumereq;
  assign _T_1287 = _T_1285 & _T_1286;
  assign haltedStatus_0 = {{31'd0}, haltedBitRegs_0};
  assign haltedSummary = haltedStatus_0 != 32'h0;
  assign _T_1323 = {{31'd0}, haltedSummary};
  assign _T_1324 = _T_1323[0];
  assign _T_1325 = _T_1323[1];
  assign _T_1326 = _T_1323[2];
  assign _T_1327 = _T_1323[3];
  assign _T_1328 = _T_1323[4];
  assign _T_1329 = _T_1323[5];
  assign _T_1330 = _T_1323[6];
  assign _T_1331 = _T_1323[7];
  assign _T_1332 = _T_1323[8];
  assign _T_1333 = _T_1323[9];
  assign _T_1334 = _T_1323[10];
  assign _T_1335 = _T_1323[11];
  assign _T_1336 = _T_1323[12];
  assign _T_1337 = _T_1323[13];
  assign _T_1338 = _T_1323[14];
  assign _T_1339 = _T_1323[15];
  assign _T_1340 = _T_1323[16];
  assign _T_1341 = _T_1323[17];
  assign _T_1342 = _T_1323[18];
  assign _T_1343 = _T_1323[19];
  assign _T_1344 = _T_1323[20];
  assign _T_1345 = _T_1323[21];
  assign _T_1346 = _T_1323[22];
  assign _T_1347 = _T_1323[23];
  assign _T_1348 = _T_1323[24];
  assign _T_1349 = _T_1323[25];
  assign _T_1350 = _T_1323[26];
  assign _T_1351 = _T_1323[27];
  assign _T_1352 = _T_1323[28];
  assign _T_1353 = _T_1323[29];
  assign _T_1354 = _T_1323[30];
  assign _T_1355 = _T_1323[31];
  assign _T_1382 = _GEN_97[10:8];
  assign ABSTRACTCSWrEn = _T_5158 & _T_103513;
  assign _T_1403 = ~ io_dmactive;
  assign _GEN_23 = _T_1403 ? 3'h0 : ABSTRACTCSReg_reserved0;
  assign _GEN_24 = _T_1403 ? 5'h10 : ABSTRACTCSReg_progsize;
  assign _GEN_25 = _T_1403 ? 11'h0 : ABSTRACTCSReg_reserved1;
  assign _GEN_27 = _T_1403 ? 1'h0 : ABSTRACTCSReg_reserved2;
  assign _GEN_28 = _T_1403 ? 3'h0 : ABSTRACTCSReg_cmderr;
  assign _GEN_29 = _T_1403 ? 3'h0 : ABSTRACTCSReg_reserved3;
  assign _GEN_30 = _T_1403 ? 5'h1 : ABSTRACTCSReg_datacount;
  assign _T_1405 = _T_1403 == 1'h0;
  assign _GEN_31 = _T_103535 ? 3'h1 : _GEN_28;
  assign _T_1408 = _T_103535 == 1'h0;
  assign _T_1409 = _T_1408 & _GEN_5668;
  assign _GEN_32 = _T_1409 ? 3'h3 : _GEN_31;
  assign _T_1414 = _GEN_5668 == 1'h0;
  assign _T_1415 = _T_1408 & _T_1414;
  assign _T_1416 = _T_1415 & _GEN_5660;
  assign _GEN_33 = _T_1416 ? 3'h2 : _GEN_32;
  assign _T_1424 = _GEN_5660 == 1'h0;
  assign _T_1425 = _T_1415 & _T_1424;
  assign _T_1426 = _T_1425 & _GEN_5662;
  assign _GEN_34 = _T_1426 ? 3'h4 : _GEN_33;
  assign _T_1437 = _GEN_5662 == 1'h0;
  assign _T_1438 = _T_1425 & _T_1437;
  assign _T_1439 = ~ _T_1382;
  assign _T_1440 = ABSTRACTCSReg_cmderr & _T_1439;
  assign _GEN_35 = ABSTRACTCSWrEn ? _T_1440 : _GEN_34;
  assign _GEN_36 = _T_1438 ? _GEN_35 : _GEN_34;
  assign _GEN_37 = _T_1405 ? _GEN_36 : _GEN_28;
  assign _T_1460 = _GEN_64[11:0];
  assign _T_1462 = _GEN_64[31:16];
  assign ABSTRACTAUTOWrEn = _T_3758 & _T_103517;
  assign _GEN_38 = _T_1403 ? 16'h0 : ABSTRACTAUTOReg_autoexecprogbuf;
  assign _GEN_39 = _T_1403 ? 4'h0 : ABSTRACTAUTOReg_reserved0;
  assign _GEN_40 = _T_1403 ? 12'h0 : ABSTRACTAUTOReg_autoexecdata;
  assign _T_1473 = _T_1405 & ABSTRACTAUTOWrEn;
  assign _T_1477 = _T_1460 & 12'h1;
  assign _GEN_41 = _T_1473 ? _T_1462 : _GEN_38;
  assign _GEN_42 = _T_1473 ? _T_1477 : _GEN_40;
  assign _T_1519 = _T_6278 | _T_6274;
  assign _T_1520 = _T_6318 | _T_6314;
  assign _T_1521 = _T_6358 | _T_6354;
  assign _T_1522 = _T_6398 | _T_6394;
  assign _T_1984 = _T_4598 | _T_4594;
  assign _T_1985 = _T_4638 | _T_4634;
  assign _T_1986 = _T_4678 | _T_4674;
  assign _T_1987 = _T_4718 | _T_4714;
  assign _T_1988 = _T_4278 | _T_4274;
  assign _T_1989 = _T_4318 | _T_4314;
  assign _T_1990 = _T_4358 | _T_4354;
  assign _T_1991 = _T_4398 | _T_4394;
  assign _T_1992 = _T_4758 | _T_4754;
  assign _T_1993 = _T_4798 | _T_4794;
  assign _T_1994 = _T_4838 | _T_4834;
  assign _T_1995 = _T_4878 | _T_4874;
  assign _T_1996 = _T_5518 | _T_5514;
  assign _T_1997 = _T_5558 | _T_5554;
  assign _T_1998 = _T_5598 | _T_5594;
  assign _T_1999 = _T_5638 | _T_5634;
  assign _T_2000 = _T_6078 | _T_6074;
  assign _T_2001 = _T_6118 | _T_6114;
  assign _T_2002 = _T_6158 | _T_6154;
  assign _T_2003 = _T_6198 | _T_6194;
  assign _T_2004 = _T_3798 | _T_3794;
  assign _T_2005 = _T_3838 | _T_3834;
  assign _T_2006 = _T_3878 | _T_3874;
  assign _T_2007 = _T_3918 | _T_3914;
  assign _T_2008 = _T_4118 | _T_4114;
  assign _T_2009 = _T_4158 | _T_4154;
  assign _T_2010 = _T_4198 | _T_4194;
  assign _T_2011 = _T_4238 | _T_4234;
  assign _T_2012 = _T_5358 | _T_5354;
  assign _T_2013 = _T_5398 | _T_5394;
  assign _T_2014 = _T_5438 | _T_5434;
  assign _T_2015 = _T_5478 | _T_5474;
  assign _T_2016 = _T_5878 | _T_5874;
  assign _T_2017 = _T_5918 | _T_5914;
  assign _T_2018 = _T_5958 | _T_5954;
  assign _T_2019 = _T_5998 | _T_5994;
  assign _T_2020 = _T_4438 | _T_4434;
  assign _T_2021 = _T_4478 | _T_4474;
  assign _T_2022 = _T_4518 | _T_4514;
  assign _T_2023 = _T_4558 | _T_4554;
  assign _T_2024 = _T_3598 | _T_3594;
  assign _T_2025 = _T_3638 | _T_3634;
  assign _T_2026 = _T_3678 | _T_3674;
  assign _T_2027 = _T_3718 | _T_3714;
  assign _T_2028 = _T_5718 | _T_5714;
  assign _T_2029 = _T_5758 | _T_5754;
  assign _T_2030 = _T_5798 | _T_5794;
  assign _T_2031 = _T_5838 | _T_5834;
  assign _T_2032 = _T_5198 | _T_5194;
  assign _T_2033 = _T_5238 | _T_5234;
  assign _T_2034 = _T_5278 | _T_5274;
  assign _T_2035 = _T_5318 | _T_5314;
  assign _T_2036 = _T_4918 | _T_4914;
  assign _T_2037 = _T_4958 | _T_4954;
  assign _T_2038 = _T_4998 | _T_4994;
  assign _T_2039 = _T_5038 | _T_5034;
  assign _T_2040 = _T_3958 | _T_3954;
  assign _T_2041 = _T_3998 | _T_3994;
  assign _T_2042 = _T_4038 | _T_4034;
  assign _T_2043 = _T_4078 | _T_4074;
  assign _T_2044 = _T_6438 | _T_6434;
  assign _T_2045 = _T_6478 | _T_6474;
  assign _T_2046 = _T_6518 | _T_6514;
  assign _T_2047 = _T_6558 | _T_6554;
  assign _T_2048 = _T_1519 | _T_1520;
  assign _T_2049 = _T_2048 | _T_1521;
  assign dmiAbstractDataAccess = _T_2049 | _T_1522;
  assign _T_2050 = _T_1984 | _T_1985;
  assign _T_2051 = _T_2050 | _T_1986;
  assign _T_2052 = _T_2051 | _T_1987;
  assign _T_2053 = _T_2052 | _T_1988;
  assign _T_2054 = _T_2053 | _T_1989;
  assign _T_2055 = _T_2054 | _T_1990;
  assign _T_2056 = _T_2055 | _T_1991;
  assign _T_2057 = _T_2056 | _T_1992;
  assign _T_2058 = _T_2057 | _T_1993;
  assign _T_2059 = _T_2058 | _T_1994;
  assign _T_2060 = _T_2059 | _T_1995;
  assign _T_2061 = _T_2060 | _T_1996;
  assign _T_2062 = _T_2061 | _T_1997;
  assign _T_2063 = _T_2062 | _T_1998;
  assign _T_2064 = _T_2063 | _T_1999;
  assign _T_2065 = _T_2064 | _T_2000;
  assign _T_2066 = _T_2065 | _T_2001;
  assign _T_2067 = _T_2066 | _T_2002;
  assign _T_2068 = _T_2067 | _T_2003;
  assign _T_2069 = _T_2068 | _T_2004;
  assign _T_2070 = _T_2069 | _T_2005;
  assign _T_2071 = _T_2070 | _T_2006;
  assign _T_2072 = _T_2071 | _T_2007;
  assign _T_2073 = _T_2072 | _T_2008;
  assign _T_2074 = _T_2073 | _T_2009;
  assign _T_2075 = _T_2074 | _T_2010;
  assign _T_2076 = _T_2075 | _T_2011;
  assign _T_2077 = _T_2076 | _T_2012;
  assign _T_2078 = _T_2077 | _T_2013;
  assign _T_2079 = _T_2078 | _T_2014;
  assign _T_2080 = _T_2079 | _T_2015;
  assign _T_2081 = _T_2080 | _T_2016;
  assign _T_2082 = _T_2081 | _T_2017;
  assign _T_2083 = _T_2082 | _T_2018;
  assign _T_2084 = _T_2083 | _T_2019;
  assign _T_2085 = _T_2084 | _T_2020;
  assign _T_2086 = _T_2085 | _T_2021;
  assign _T_2087 = _T_2086 | _T_2022;
  assign _T_2088 = _T_2087 | _T_2023;
  assign _T_2089 = _T_2088 | _T_2024;
  assign _T_2090 = _T_2089 | _T_2025;
  assign _T_2091 = _T_2090 | _T_2026;
  assign _T_2092 = _T_2091 | _T_2027;
  assign _T_2093 = _T_2092 | _T_2028;
  assign _T_2094 = _T_2093 | _T_2029;
  assign _T_2095 = _T_2094 | _T_2030;
  assign _T_2096 = _T_2095 | _T_2031;
  assign _T_2097 = _T_2096 | _T_2032;
  assign _T_2098 = _T_2097 | _T_2033;
  assign _T_2099 = _T_2098 | _T_2034;
  assign _T_2100 = _T_2099 | _T_2035;
  assign _T_2101 = _T_2100 | _T_2036;
  assign _T_2102 = _T_2101 | _T_2037;
  assign _T_2103 = _T_2102 | _T_2038;
  assign _T_2104 = _T_2103 | _T_2039;
  assign _T_2105 = _T_2104 | _T_2040;
  assign _T_2106 = _T_2105 | _T_2041;
  assign _T_2107 = _T_2106 | _T_2042;
  assign _T_2108 = _T_2107 | _T_2043;
  assign _T_2109 = _T_2108 | _T_2044;
  assign _T_2110 = _T_2109 | _T_2045;
  assign _T_2111 = _T_2110 | _T_2046;
  assign dmiProgramBufferAccess = _T_2111 | _T_2047;
  assign _T_2257 = ABSTRACTAUTOReg_autoexecdata[0];
  assign _T_2269 = _T_1519 & _T_2257;
  assign _T_2270 = ABSTRACTAUTOReg_autoexecprogbuf[0];
  assign _T_2271 = ABSTRACTAUTOReg_autoexecprogbuf[1];
  assign _T_2272 = ABSTRACTAUTOReg_autoexecprogbuf[2];
  assign _T_2273 = ABSTRACTAUTOReg_autoexecprogbuf[3];
  assign _T_2274 = ABSTRACTAUTOReg_autoexecprogbuf[4];
  assign _T_2275 = ABSTRACTAUTOReg_autoexecprogbuf[5];
  assign _T_2276 = ABSTRACTAUTOReg_autoexecprogbuf[6];
  assign _T_2277 = ABSTRACTAUTOReg_autoexecprogbuf[7];
  assign _T_2278 = ABSTRACTAUTOReg_autoexecprogbuf[8];
  assign _T_2279 = ABSTRACTAUTOReg_autoexecprogbuf[9];
  assign _T_2280 = ABSTRACTAUTOReg_autoexecprogbuf[10];
  assign _T_2281 = ABSTRACTAUTOReg_autoexecprogbuf[11];
  assign _T_2282 = ABSTRACTAUTOReg_autoexecprogbuf[12];
  assign _T_2283 = ABSTRACTAUTOReg_autoexecprogbuf[13];
  assign _T_2284 = ABSTRACTAUTOReg_autoexecprogbuf[14];
  assign _T_2285 = ABSTRACTAUTOReg_autoexecprogbuf[15];
  assign _T_2286 = _T_1984 & _T_2270;
  assign _T_2287 = _T_1988 & _T_2271;
  assign _T_2288 = _T_1992 & _T_2272;
  assign _T_2289 = _T_1996 & _T_2273;
  assign _T_2290 = _T_2000 & _T_2274;
  assign _T_2291 = _T_2004 & _T_2275;
  assign _T_2292 = _T_2008 & _T_2276;
  assign _T_2293 = _T_2012 & _T_2277;
  assign _T_2294 = _T_2016 & _T_2278;
  assign _T_2295 = _T_2020 & _T_2279;
  assign _T_2296 = _T_2024 & _T_2280;
  assign _T_2297 = _T_2028 & _T_2281;
  assign _T_2298 = _T_2032 & _T_2282;
  assign _T_2299 = _T_2036 & _T_2283;
  assign _T_2300 = _T_2040 & _T_2284;
  assign _T_2301 = _T_2044 & _T_2285;
  assign _T_2302 = _T_2286 | _T_2287;
  assign _T_2303 = _T_2302 | _T_2288;
  assign _T_2304 = _T_2303 | _T_2289;
  assign _T_2305 = _T_2304 | _T_2290;
  assign _T_2306 = _T_2305 | _T_2291;
  assign _T_2307 = _T_2306 | _T_2292;
  assign _T_2308 = _T_2307 | _T_2293;
  assign _T_2309 = _T_2308 | _T_2294;
  assign _T_2310 = _T_2309 | _T_2295;
  assign _T_2311 = _T_2310 | _T_2296;
  assign _T_2312 = _T_2311 | _T_2297;
  assign _T_2313 = _T_2312 | _T_2298;
  assign _T_2314 = _T_2313 | _T_2299;
  assign _T_2315 = _T_2314 | _T_2300;
  assign _T_2316 = _T_2315 | _T_2301;
  assign autoexec = _T_2269 | _T_2316;
  assign _T_2334 = _GEN_118[23:0];
  assign _T_2335 = _GEN_118[31:24];
  assign COMMANDWrEn = _T_6038 & _T_103515;
  assign _GEN_43 = _T_1403 ? 8'h0 : COMMANDRdData_cmdtype;
  assign _GEN_44 = _T_1403 ? 24'h0 : COMMANDRdData_control;
  assign _GEN_45 = COMMANDWrEn ? _T_2335 : _GEN_43;
  assign _GEN_46 = COMMANDWrEn ? _T_2334 : _GEN_44;
  assign _GEN_47 = _T_1405 ? _GEN_45 : _GEN_43;
  assign _GEN_48 = _T_1405 ? _GEN_46 : _GEN_44;
  assign _GEN_49 = _T_1403 ? 1'h0 : haltedBitRegs_0;
  assign _GEN_50 = _T_1403 ? 1'h0 : resumeReqRegs_0;
  assign _T_2786 = _T_57264 == 10'h0;
  assign _GEN_51 = _T_2786 ? 1'h1 : _GEN_49;
  assign _GEN_52 = _T_57263 ? _GEN_51 : _GEN_49;
  assign _T_2789 = _T_57263 == 1'h0;
  assign _T_2790 = _T_2789 & _T_63863;
  assign _T_2792 = _T_63864 == 10'h0;
  assign _GEN_53 = _T_2792 ? 1'h0 : _GEN_52;
  assign _GEN_54 = _T_2790 ? _GEN_53 : _GEN_52;
  assign _GEN_55 = _T_2792 ? 1'h0 : _GEN_50;
  assign _GEN_56 = _T_63863 ? _GEN_55 : _GEN_50;
  assign _GEN_57 = resumereq ? 1'h1 : _GEN_56;
  assign _GEN_58 = _T_1405 ? _GEN_54 : _GEN_49;
  assign _GEN_59 = _T_1405 ? _GEN_57 : _GEN_50;
  assign _T_2806 = {_T_1267,_T_1267};
  assign _T_2807 = {_T_2806,2'h2};
  assign _T_2808 = {_T_2807,6'h2};
  assign _T_2809 = {_T_1277,_T_1277};
  assign _T_2810 = {_T_1255,_T_1255};
  assign _T_2811 = {_T_2810,_T_2809};
  assign _T_2812 = {_T_1246,_T_1246};
  assign _T_2813 = {14'h0,_T_1287};
  assign _T_2814 = {_T_2813,_T_1287};
  assign _T_2815 = {_T_2814,_T_2812};
  assign _T_2816 = {_T_2815,_T_2811};
  assign _T_2817 = {_T_2816,_T_2808};
  assign _T_2823 = {_T_1325,_T_1324};
  assign _T_2824 = {_T_1327,_T_1326};
  assign _T_2825 = {_T_2824,_T_2823};
  assign _T_2826 = {_T_1329,_T_1328};
  assign _T_2827 = {_T_1331,_T_1330};
  assign _T_2828 = {_T_2827,_T_2826};
  assign _T_2829 = {_T_2828,_T_2825};
  assign _T_2830 = {_T_1333,_T_1332};
  assign _T_2831 = {_T_1335,_T_1334};
  assign _T_2832 = {_T_2831,_T_2830};
  assign _T_2833 = {_T_1337,_T_1336};
  assign _T_2834 = {_T_1339,_T_1338};
  assign _T_2835 = {_T_2834,_T_2833};
  assign _T_2836 = {_T_2835,_T_2832};
  assign _T_2837 = {_T_2836,_T_2829};
  assign _T_2838 = {_T_1341,_T_1340};
  assign _T_2839 = {_T_1343,_T_1342};
  assign _T_2840 = {_T_2839,_T_2838};
  assign _T_2841 = {_T_1345,_T_1344};
  assign _T_2842 = {_T_1347,_T_1346};
  assign _T_2843 = {_T_2842,_T_2841};
  assign _T_2844 = {_T_2843,_T_2840};
  assign _T_2845 = {_T_1349,_T_1348};
  assign _T_2846 = {_T_1351,_T_1350};
  assign _T_2847 = {_T_2846,_T_2845};
  assign _T_2848 = {_T_1353,_T_1352};
  assign _T_2849 = {_T_1355,_T_1354};
  assign _T_2850 = {_T_2849,_T_2848};
  assign _T_2851 = {_T_2850,_T_2847};
  assign _T_2852 = {_T_2851,_T_2844};
  assign _T_2853 = {_T_2852,_T_2837};
  assign _T_2854 = {ABSTRACTCSReg_reserved3,ABSTRACTCSReg_datacount};
  assign _T_2855 = {ABSTRACTCSReg_reserved2,ABSTRACTCSReg_cmderr};
  assign _T_2856 = {_T_2855,_T_2854};
  assign _T_2857 = {ABSTRACTCSReg_reserved1,_T_103511};
  assign _T_2858 = {ABSTRACTCSReg_reserved0,ABSTRACTCSReg_progsize};
  assign _T_2859 = {_T_2858,_T_2857};
  assign _T_2860 = {_T_2859,_T_2856};
  assign _T_2861 = {ABSTRACTAUTOReg_autoexecprogbuf,ABSTRACTAUTOReg_reserved0};
  assign _T_2862 = {_T_2861,ABSTRACTAUTOReg_autoexecdata};
  assign _T_2863 = {COMMANDRdData_cmdtype,COMMANDRdData_control};
  assign _T_2874 = io_dmi_in_0_a_bits_opcode == 3'h4;
  assign _T_2875 = io_dmi_in_0_a_bits_address[8:2];
  assign _T_2876 = {io_dmi_in_0_a_bits_source,io_dmi_in_0_a_bits_size};
  assign _T_2962 = _T_2875 ^ 7'h2a;
  assign _T_2963 = _T_2962 & 7'h50;
  assign _T_2965 = _T_2963 == 7'h0;
  assign _T_2971 = _T_2875 ^ 7'h18;
  assign _T_2972 = _T_2971 & 7'h50;
  assign _T_2974 = _T_2972 == 7'h0;
  assign _T_2980 = _T_2875 ^ 7'h25;
  assign _T_2981 = _T_2980 & 7'h50;
  assign _T_2983 = _T_2981 == 7'h0;
  assign _T_2989 = _T_2875 ^ 7'h2e;
  assign _T_2990 = _T_2989 & 7'h50;
  assign _T_2992 = _T_2990 == 7'h0;
  assign _T_2998 = _T_2875 ^ 7'h26;
  assign _T_2999 = _T_2998 & 7'h50;
  assign _T_3001 = _T_2999 == 7'h0;
  assign _T_3007 = _T_2875 ^ 7'h21;
  assign _T_3008 = _T_3007 & 7'h50;
  assign _T_3010 = _T_3008 == 7'h0;
  assign _T_3016 = _T_2875 ^ 7'h29;
  assign _T_3017 = _T_3016 & 7'h50;
  assign _T_3019 = _T_3017 == 7'h0;
  assign _T_3025 = _T_2875 ^ 7'h20;
  assign _T_3026 = _T_3025 & 7'h50;
  assign _T_3028 = _T_3026 == 7'h0;
  assign _T_3034 = _T_2875 ^ 7'h22;
  assign _T_3035 = _T_3034 & 7'h50;
  assign _T_3037 = _T_3035 == 7'h0;
  assign _T_3043 = _T_2875 ^ 7'h2d;
  assign _T_3044 = _T_3043 & 7'h50;
  assign _T_3046 = _T_3044 == 7'h0;
  assign _T_3052 = _T_2875 ^ 7'h40;
  assign _T_3053 = _T_3052 & 7'h50;
  assign _T_3055 = _T_3053 == 7'h0;
  assign _T_3061 = _T_2875 ^ 7'h11;
  assign _T_3062 = _T_3061 & 7'h50;
  assign _T_3064 = _T_3062 == 7'h0;
  assign _T_3070 = _T_2875 ^ 7'h16;
  assign _T_3071 = _T_3070 & 7'h50;
  assign _T_3073 = _T_3071 == 7'h0;
  assign _T_3079 = _T_2875 ^ 7'h2c;
  assign _T_3080 = _T_3079 & 7'h50;
  assign _T_3082 = _T_3080 == 7'h0;
  assign _T_3088 = _T_2875 ^ 7'h27;
  assign _T_3089 = _T_3088 & 7'h50;
  assign _T_3091 = _T_3089 == 7'h0;
  assign _T_3097 = _T_2875 ^ 7'h23;
  assign _T_3098 = _T_3097 & 7'h50;
  assign _T_3100 = _T_3098 == 7'h0;
  assign _T_3106 = _T_2875 ^ 7'h12;
  assign _T_3107 = _T_3106 & 7'h50;
  assign _T_3109 = _T_3107 == 7'h0;
  assign _T_3115 = _T_2875 ^ 7'h2b;
  assign _T_3116 = _T_3115 & 7'h50;
  assign _T_3118 = _T_3116 == 7'h0;
  assign _T_3124 = _T_2875 ^ 7'h28;
  assign _T_3125 = _T_3124 & 7'h50;
  assign _T_3127 = _T_3125 == 7'h0;
  assign _T_3133 = _T_2875 ^ 7'h17;
  assign _T_3134 = _T_3133 & 7'h50;
  assign _T_3136 = _T_3134 == 7'h0;
  assign _T_3142 = _T_2875 ^ 7'h24;
  assign _T_3143 = _T_3142 & 7'h50;
  assign _T_3145 = _T_3143 == 7'h0;
  assign _T_3151 = _T_2875 ^ 7'h13;
  assign _T_3152 = _T_3151 & 7'h50;
  assign _T_3154 = _T_3152 == 7'h0;
  assign _T_3160 = _T_2875 ^ 7'h4;
  assign _T_3161 = _T_3160 & 7'h50;
  assign _T_3163 = _T_3161 == 7'h0;
  assign _T_3169 = _T_2875 ^ 7'h2f;
  assign _T_3170 = _T_3169 & 7'h50;
  assign _T_3172 = _T_3170 == 7'h0;
  assign _T_3533 = io_dmi_in_0_a_bits_mask[0];
  assign _T_3534 = io_dmi_in_0_a_bits_mask[1];
  assign _T_3535 = io_dmi_in_0_a_bits_mask[2];
  assign _T_3536 = io_dmi_in_0_a_bits_mask[3];
  assign _T_3540 = _T_3533 ? 8'hff : 8'h0;
  assign _T_3544 = _T_3534 ? 8'hff : 8'h0;
  assign _T_3548 = _T_3535 ? 8'hff : 8'h0;
  assign _T_3552 = _T_3536 ? 8'hff : 8'h0;
  assign _T_3553 = {_T_3544,_T_3540};
  assign _T_3554 = {_T_3552,_T_3548};
  assign _T_3555 = {_T_3554,_T_3553};
  assign _T_3579 = _T_3555[7:0];
  assign _T_3581 = _T_3579 != 8'h0;
  assign _T_3583 = ~ _T_3579;
  assign _T_3585 = _T_3583 == 8'h0;
  assign _T_3594 = _T_7474 & _T_3581;
  assign _T_3598 = _T_7771 & _T_3585;
  assign _T_3599 = io_dmi_in_0_a_bits_data[7:0];
  assign _GEN_60 = _T_3598 ? _T_3599 : programBufferMem_40;
  assign _T_3619 = _T_3555[15:8];
  assign _T_3621 = _T_3619 != 8'h0;
  assign _T_3623 = ~ _T_3619;
  assign _T_3625 = _T_3623 == 8'h0;
  assign _T_3634 = _T_7474 & _T_3621;
  assign _T_3638 = _T_7771 & _T_3625;
  assign _T_3639 = io_dmi_in_0_a_bits_data[15:8];
  assign _GEN_61 = _T_3638 ? _T_3639 : programBufferMem_41;
  assign _GEN_5671 = {{8'd0}, programBufferMem_41};
  assign _T_3654 = _GEN_5671 << 8;
  assign _GEN_5672 = {{8'd0}, programBufferMem_40};
  assign _T_3658 = _GEN_5672 | _T_3654;
  assign _T_3659 = _T_3555[23:16];
  assign _T_3661 = _T_3659 != 8'h0;
  assign _T_3663 = ~ _T_3659;
  assign _T_3665 = _T_3663 == 8'h0;
  assign _T_3674 = _T_7474 & _T_3661;
  assign _T_3678 = _T_7771 & _T_3665;
  assign _T_3679 = io_dmi_in_0_a_bits_data[23:16];
  assign _GEN_62 = _T_3678 ? _T_3679 : programBufferMem_42;
  assign _GEN_5673 = {{16'd0}, programBufferMem_42};
  assign _T_3694 = _GEN_5673 << 16;
  assign _GEN_5674 = {{8'd0}, _T_3658};
  assign _T_3698 = _GEN_5674 | _T_3694;
  assign _T_3699 = _T_3555[31:24];
  assign _T_3701 = _T_3699 != 8'h0;
  assign _T_3703 = ~ _T_3699;
  assign _T_3705 = _T_3703 == 8'h0;
  assign _T_3714 = _T_7474 & _T_3701;
  assign _T_3718 = _T_7771 & _T_3705;
  assign _T_3719 = io_dmi_in_0_a_bits_data[31:24];
  assign _GEN_63 = _T_3718 ? _T_3719 : programBufferMem_43;
  assign _GEN_5675 = {{24'd0}, programBufferMem_43};
  assign _T_3734 = _GEN_5675 << 24;
  assign _GEN_5676 = {{8'd0}, _T_3698};
  assign _T_3738 = _GEN_5676 | _T_3734;
  assign _T_3743 = ~ _T_3555;
  assign _T_3745 = _T_3743 == 32'h0;
  assign _T_3758 = _T_7627 & _T_3745;
  assign _GEN_64 = _T_3758 ? io_dmi_in_0_a_bits_data : 32'h0;
  assign _T_3794 = _T_7434 & _T_3581;
  assign _T_3798 = _T_7731 & _T_3585;
  assign _GEN_65 = _T_3798 ? _T_3599 : programBufferMem_20;
  assign _T_3834 = _T_7434 & _T_3621;
  assign _T_3838 = _T_7731 & _T_3625;
  assign _GEN_66 = _T_3838 ? _T_3639 : programBufferMem_21;
  assign _GEN_5677 = {{8'd0}, programBufferMem_21};
  assign _T_3854 = _GEN_5677 << 8;
  assign _GEN_5678 = {{8'd0}, programBufferMem_20};
  assign _T_3858 = _GEN_5678 | _T_3854;
  assign _T_3874 = _T_7434 & _T_3661;
  assign _T_3878 = _T_7731 & _T_3665;
  assign _GEN_67 = _T_3878 ? _T_3679 : programBufferMem_22;
  assign _GEN_5679 = {{16'd0}, programBufferMem_22};
  assign _T_3894 = _GEN_5679 << 16;
  assign _GEN_5680 = {{8'd0}, _T_3858};
  assign _T_3898 = _GEN_5680 | _T_3894;
  assign _T_3914 = _T_7434 & _T_3701;
  assign _T_3918 = _T_7731 & _T_3705;
  assign _GEN_68 = _T_3918 ? _T_3719 : programBufferMem_23;
  assign _GEN_5681 = {{24'd0}, programBufferMem_23};
  assign _T_3934 = _GEN_5681 << 24;
  assign _GEN_5682 = {{8'd0}, _T_3898};
  assign _T_3938 = _GEN_5682 | _T_3934;
  assign _T_3954 = _T_7506 & _T_3581;
  assign _T_3958 = _T_7803 & _T_3585;
  assign _GEN_69 = _T_3958 ? _T_3599 : programBufferMem_56;
  assign _T_3994 = _T_7506 & _T_3621;
  assign _T_3998 = _T_7803 & _T_3625;
  assign _GEN_70 = _T_3998 ? _T_3639 : programBufferMem_57;
  assign _GEN_5683 = {{8'd0}, programBufferMem_57};
  assign _T_4014 = _GEN_5683 << 8;
  assign _GEN_5684 = {{8'd0}, programBufferMem_56};
  assign _T_4018 = _GEN_5684 | _T_4014;
  assign _T_4034 = _T_7506 & _T_3661;
  assign _T_4038 = _T_7803 & _T_3665;
  assign _GEN_71 = _T_4038 ? _T_3679 : programBufferMem_58;
  assign _GEN_5685 = {{16'd0}, programBufferMem_58};
  assign _T_4054 = _GEN_5685 << 16;
  assign _GEN_5686 = {{8'd0}, _T_4018};
  assign _T_4058 = _GEN_5686 | _T_4054;
  assign _T_4074 = _T_7506 & _T_3701;
  assign _T_4078 = _T_7803 & _T_3705;
  assign _GEN_72 = _T_4078 ? _T_3719 : programBufferMem_59;
  assign _GEN_5687 = {{24'd0}, programBufferMem_59};
  assign _T_4094 = _GEN_5687 << 24;
  assign _GEN_5688 = {{8'd0}, _T_4058};
  assign _T_4098 = _GEN_5688 | _T_4094;
  assign _T_4114 = _T_7442 & _T_3581;
  assign _T_4118 = _T_7739 & _T_3585;
  assign _GEN_73 = _T_4118 ? _T_3599 : programBufferMem_24;
  assign _T_4154 = _T_7442 & _T_3621;
  assign _T_4158 = _T_7739 & _T_3625;
  assign _GEN_74 = _T_4158 ? _T_3639 : programBufferMem_25;
  assign _GEN_5689 = {{8'd0}, programBufferMem_25};
  assign _T_4174 = _GEN_5689 << 8;
  assign _GEN_5690 = {{8'd0}, programBufferMem_24};
  assign _T_4178 = _GEN_5690 | _T_4174;
  assign _T_4194 = _T_7442 & _T_3661;
  assign _T_4198 = _T_7739 & _T_3665;
  assign _GEN_75 = _T_4198 ? _T_3679 : programBufferMem_26;
  assign _GEN_5691 = {{16'd0}, programBufferMem_26};
  assign _T_4214 = _GEN_5691 << 16;
  assign _GEN_5692 = {{8'd0}, _T_4178};
  assign _T_4218 = _GEN_5692 | _T_4214;
  assign _T_4234 = _T_7442 & _T_3701;
  assign _T_4238 = _T_7739 & _T_3705;
  assign _GEN_76 = _T_4238 ? _T_3719 : programBufferMem_27;
  assign _GEN_5693 = {{24'd0}, programBufferMem_27};
  assign _T_4254 = _GEN_5693 << 24;
  assign _GEN_5694 = {{8'd0}, _T_4218};
  assign _T_4258 = _GEN_5694 | _T_4254;
  assign _T_4274 = _T_7402 & _T_3581;
  assign _T_4278 = _T_7699 & _T_3585;
  assign _GEN_77 = _T_4278 ? _T_3599 : programBufferMem_4;
  assign _T_4314 = _T_7402 & _T_3621;
  assign _T_4318 = _T_7699 & _T_3625;
  assign _GEN_78 = _T_4318 ? _T_3639 : programBufferMem_5;
  assign _GEN_5695 = {{8'd0}, programBufferMem_5};
  assign _T_4334 = _GEN_5695 << 8;
  assign _GEN_5696 = {{8'd0}, programBufferMem_4};
  assign _T_4338 = _GEN_5696 | _T_4334;
  assign _T_4354 = _T_7402 & _T_3661;
  assign _T_4358 = _T_7699 & _T_3665;
  assign _GEN_79 = _T_4358 ? _T_3679 : programBufferMem_6;
  assign _GEN_5697 = {{16'd0}, programBufferMem_6};
  assign _T_4374 = _GEN_5697 << 16;
  assign _GEN_5698 = {{8'd0}, _T_4338};
  assign _T_4378 = _GEN_5698 | _T_4374;
  assign _T_4394 = _T_7402 & _T_3701;
  assign _T_4398 = _T_7699 & _T_3705;
  assign _GEN_80 = _T_4398 ? _T_3719 : programBufferMem_7;
  assign _GEN_5699 = {{24'd0}, programBufferMem_7};
  assign _T_4414 = _GEN_5699 << 24;
  assign _GEN_5700 = {{8'd0}, _T_4378};
  assign _T_4418 = _GEN_5700 | _T_4414;
  assign _T_4434 = _T_7466 & _T_3581;
  assign _T_4438 = _T_7763 & _T_3585;
  assign _GEN_81 = _T_4438 ? _T_3599 : programBufferMem_36;
  assign _T_4474 = _T_7466 & _T_3621;
  assign _T_4478 = _T_7763 & _T_3625;
  assign _GEN_82 = _T_4478 ? _T_3639 : programBufferMem_37;
  assign _GEN_5701 = {{8'd0}, programBufferMem_37};
  assign _T_4494 = _GEN_5701 << 8;
  assign _GEN_5702 = {{8'd0}, programBufferMem_36};
  assign _T_4498 = _GEN_5702 | _T_4494;
  assign _T_4514 = _T_7466 & _T_3661;
  assign _T_4518 = _T_7763 & _T_3665;
  assign _GEN_83 = _T_4518 ? _T_3679 : programBufferMem_38;
  assign _GEN_5703 = {{16'd0}, programBufferMem_38};
  assign _T_4534 = _GEN_5703 << 16;
  assign _GEN_5704 = {{8'd0}, _T_4498};
  assign _T_4538 = _GEN_5704 | _T_4534;
  assign _T_4554 = _T_7466 & _T_3701;
  assign _T_4558 = _T_7763 & _T_3705;
  assign _GEN_84 = _T_4558 ? _T_3719 : programBufferMem_39;
  assign _GEN_5705 = {{24'd0}, programBufferMem_39};
  assign _T_4574 = _GEN_5705 << 24;
  assign _GEN_5706 = {{8'd0}, _T_4538};
  assign _T_4578 = _GEN_5706 | _T_4574;
  assign _T_4594 = _T_7394 & _T_3581;
  assign _T_4598 = _T_7691 & _T_3585;
  assign _GEN_85 = _T_4598 ? _T_3599 : programBufferMem_0;
  assign _T_4634 = _T_7394 & _T_3621;
  assign _T_4638 = _T_7691 & _T_3625;
  assign _GEN_86 = _T_4638 ? _T_3639 : programBufferMem_1;
  assign _GEN_5707 = {{8'd0}, programBufferMem_1};
  assign _T_4654 = _GEN_5707 << 8;
  assign _GEN_5708 = {{8'd0}, programBufferMem_0};
  assign _T_4658 = _GEN_5708 | _T_4654;
  assign _T_4674 = _T_7394 & _T_3661;
  assign _T_4678 = _T_7691 & _T_3665;
  assign _GEN_87 = _T_4678 ? _T_3679 : programBufferMem_2;
  assign _GEN_5709 = {{16'd0}, programBufferMem_2};
  assign _T_4694 = _GEN_5709 << 16;
  assign _GEN_5710 = {{8'd0}, _T_4658};
  assign _T_4698 = _GEN_5710 | _T_4694;
  assign _T_4714 = _T_7394 & _T_3701;
  assign _T_4718 = _T_7691 & _T_3705;
  assign _GEN_88 = _T_4718 ? _T_3719 : programBufferMem_3;
  assign _GEN_5711 = {{24'd0}, programBufferMem_3};
  assign _T_4734 = _GEN_5711 << 24;
  assign _GEN_5712 = {{8'd0}, _T_4698};
  assign _T_4738 = _GEN_5712 | _T_4734;
  assign _T_4754 = _T_7410 & _T_3581;
  assign _T_4758 = _T_7707 & _T_3585;
  assign _GEN_89 = _T_4758 ? _T_3599 : programBufferMem_8;
  assign _T_4794 = _T_7410 & _T_3621;
  assign _T_4798 = _T_7707 & _T_3625;
  assign _GEN_90 = _T_4798 ? _T_3639 : programBufferMem_9;
  assign _GEN_5713 = {{8'd0}, programBufferMem_9};
  assign _T_4814 = _GEN_5713 << 8;
  assign _GEN_5714 = {{8'd0}, programBufferMem_8};
  assign _T_4818 = _GEN_5714 | _T_4814;
  assign _T_4834 = _T_7410 & _T_3661;
  assign _T_4838 = _T_7707 & _T_3665;
  assign _GEN_91 = _T_4838 ? _T_3679 : programBufferMem_10;
  assign _GEN_5715 = {{16'd0}, programBufferMem_10};
  assign _T_4854 = _GEN_5715 << 16;
  assign _GEN_5716 = {{8'd0}, _T_4818};
  assign _T_4858 = _GEN_5716 | _T_4854;
  assign _T_4874 = _T_7410 & _T_3701;
  assign _T_4878 = _T_7707 & _T_3705;
  assign _GEN_92 = _T_4878 ? _T_3719 : programBufferMem_11;
  assign _GEN_5717 = {{24'd0}, programBufferMem_11};
  assign _T_4894 = _GEN_5717 << 24;
  assign _GEN_5718 = {{8'd0}, _T_4858};
  assign _T_4898 = _GEN_5718 | _T_4894;
  assign _T_4914 = _T_7498 & _T_3581;
  assign _T_4918 = _T_7795 & _T_3585;
  assign _GEN_93 = _T_4918 ? _T_3599 : programBufferMem_52;
  assign _T_4954 = _T_7498 & _T_3621;
  assign _T_4958 = _T_7795 & _T_3625;
  assign _GEN_94 = _T_4958 ? _T_3639 : programBufferMem_53;
  assign _GEN_5719 = {{8'd0}, programBufferMem_53};
  assign _T_4974 = _GEN_5719 << 8;
  assign _GEN_5720 = {{8'd0}, programBufferMem_52};
  assign _T_4978 = _GEN_5720 | _T_4974;
  assign _T_4994 = _T_7498 & _T_3661;
  assign _T_4998 = _T_7795 & _T_3665;
  assign _GEN_95 = _T_4998 ? _T_3679 : programBufferMem_54;
  assign _GEN_5721 = {{16'd0}, programBufferMem_54};
  assign _T_5014 = _GEN_5721 << 16;
  assign _GEN_5722 = {{8'd0}, _T_4978};
  assign _T_5018 = _GEN_5722 | _T_5014;
  assign _T_5034 = _T_7498 & _T_3701;
  assign _T_5038 = _T_7795 & _T_3705;
  assign _GEN_96 = _T_5038 ? _T_3719 : programBufferMem_55;
  assign _GEN_5723 = {{24'd0}, programBufferMem_55};
  assign _T_5054 = _GEN_5723 << 24;
  assign _GEN_5724 = {{8'd0}, _T_5018};
  assign _T_5058 = _GEN_5724 | _T_5054;
  assign _T_5158 = _T_7611 & _T_3745;
  assign _GEN_97 = _T_5158 ? io_dmi_in_0_a_bits_data : 32'h0;
  assign _T_5194 = _T_7490 & _T_3581;
  assign _T_5198 = _T_7787 & _T_3585;
  assign _GEN_98 = _T_5198 ? _T_3599 : programBufferMem_48;
  assign _T_5234 = _T_7490 & _T_3621;
  assign _T_5238 = _T_7787 & _T_3625;
  assign _GEN_99 = _T_5238 ? _T_3639 : programBufferMem_49;
  assign _GEN_5725 = {{8'd0}, programBufferMem_49};
  assign _T_5254 = _GEN_5725 << 8;
  assign _GEN_5726 = {{8'd0}, programBufferMem_48};
  assign _T_5258 = _GEN_5726 | _T_5254;
  assign _T_5274 = _T_7490 & _T_3661;
  assign _T_5278 = _T_7787 & _T_3665;
  assign _GEN_100 = _T_5278 ? _T_3679 : programBufferMem_50;
  assign _GEN_5727 = {{16'd0}, programBufferMem_50};
  assign _T_5294 = _GEN_5727 << 16;
  assign _GEN_5728 = {{8'd0}, _T_5258};
  assign _T_5298 = _GEN_5728 | _T_5294;
  assign _T_5314 = _T_7490 & _T_3701;
  assign _T_5318 = _T_7787 & _T_3705;
  assign _GEN_101 = _T_5318 ? _T_3719 : programBufferMem_51;
  assign _GEN_5729 = {{24'd0}, programBufferMem_51};
  assign _T_5334 = _GEN_5729 << 24;
  assign _GEN_5730 = {{8'd0}, _T_5298};
  assign _T_5338 = _GEN_5730 | _T_5334;
  assign _T_5354 = _T_7450 & _T_3581;
  assign _T_5358 = _T_7747 & _T_3585;
  assign _GEN_102 = _T_5358 ? _T_3599 : programBufferMem_28;
  assign _T_5394 = _T_7450 & _T_3621;
  assign _T_5398 = _T_7747 & _T_3625;
  assign _GEN_103 = _T_5398 ? _T_3639 : programBufferMem_29;
  assign _GEN_5731 = {{8'd0}, programBufferMem_29};
  assign _T_5414 = _GEN_5731 << 8;
  assign _GEN_5732 = {{8'd0}, programBufferMem_28};
  assign _T_5418 = _GEN_5732 | _T_5414;
  assign _T_5434 = _T_7450 & _T_3661;
  assign _T_5438 = _T_7747 & _T_3665;
  assign _GEN_104 = _T_5438 ? _T_3679 : programBufferMem_30;
  assign _GEN_5733 = {{16'd0}, programBufferMem_30};
  assign _T_5454 = _GEN_5733 << 16;
  assign _GEN_5734 = {{8'd0}, _T_5418};
  assign _T_5458 = _GEN_5734 | _T_5454;
  assign _T_5474 = _T_7450 & _T_3701;
  assign _T_5478 = _T_7747 & _T_3705;
  assign _GEN_105 = _T_5478 ? _T_3719 : programBufferMem_31;
  assign _GEN_5735 = {{24'd0}, programBufferMem_31};
  assign _T_5494 = _GEN_5735 << 24;
  assign _GEN_5736 = {{8'd0}, _T_5458};
  assign _T_5498 = _GEN_5736 | _T_5494;
  assign _T_5514 = _T_7418 & _T_3581;
  assign _T_5518 = _T_7715 & _T_3585;
  assign _GEN_106 = _T_5518 ? _T_3599 : programBufferMem_12;
  assign _T_5554 = _T_7418 & _T_3621;
  assign _T_5558 = _T_7715 & _T_3625;
  assign _GEN_107 = _T_5558 ? _T_3639 : programBufferMem_13;
  assign _GEN_5737 = {{8'd0}, programBufferMem_13};
  assign _T_5574 = _GEN_5737 << 8;
  assign _GEN_5738 = {{8'd0}, programBufferMem_12};
  assign _T_5578 = _GEN_5738 | _T_5574;
  assign _T_5594 = _T_7418 & _T_3661;
  assign _T_5598 = _T_7715 & _T_3665;
  assign _GEN_108 = _T_5598 ? _T_3679 : programBufferMem_14;
  assign _GEN_5739 = {{16'd0}, programBufferMem_14};
  assign _T_5614 = _GEN_5739 << 16;
  assign _GEN_5740 = {{8'd0}, _T_5578};
  assign _T_5618 = _GEN_5740 | _T_5614;
  assign _T_5634 = _T_7418 & _T_3701;
  assign _T_5638 = _T_7715 & _T_3705;
  assign _GEN_109 = _T_5638 ? _T_3719 : programBufferMem_15;
  assign _GEN_5741 = {{24'd0}, programBufferMem_15};
  assign _T_5654 = _GEN_5741 << 24;
  assign _GEN_5742 = {{8'd0}, _T_5618};
  assign _T_5658 = _GEN_5742 | _T_5654;
  assign _T_5714 = _T_7482 & _T_3581;
  assign _T_5718 = _T_7779 & _T_3585;
  assign _GEN_110 = _T_5718 ? _T_3599 : programBufferMem_44;
  assign _T_5754 = _T_7482 & _T_3621;
  assign _T_5758 = _T_7779 & _T_3625;
  assign _GEN_111 = _T_5758 ? _T_3639 : programBufferMem_45;
  assign _GEN_5743 = {{8'd0}, programBufferMem_45};
  assign _T_5774 = _GEN_5743 << 8;
  assign _GEN_5744 = {{8'd0}, programBufferMem_44};
  assign _T_5778 = _GEN_5744 | _T_5774;
  assign _T_5794 = _T_7482 & _T_3661;
  assign _T_5798 = _T_7779 & _T_3665;
  assign _GEN_112 = _T_5798 ? _T_3679 : programBufferMem_46;
  assign _GEN_5745 = {{16'd0}, programBufferMem_46};
  assign _T_5814 = _GEN_5745 << 16;
  assign _GEN_5746 = {{8'd0}, _T_5778};
  assign _T_5818 = _GEN_5746 | _T_5814;
  assign _T_5834 = _T_7482 & _T_3701;
  assign _T_5838 = _T_7779 & _T_3705;
  assign _GEN_113 = _T_5838 ? _T_3719 : programBufferMem_47;
  assign _GEN_5747 = {{24'd0}, programBufferMem_47};
  assign _T_5854 = _GEN_5747 << 24;
  assign _GEN_5748 = {{8'd0}, _T_5818};
  assign _T_5858 = _GEN_5748 | _T_5854;
  assign _T_5874 = _T_7458 & _T_3581;
  assign _T_5878 = _T_7755 & _T_3585;
  assign _GEN_114 = _T_5878 ? _T_3599 : programBufferMem_32;
  assign _T_5914 = _T_7458 & _T_3621;
  assign _T_5918 = _T_7755 & _T_3625;
  assign _GEN_115 = _T_5918 ? _T_3639 : programBufferMem_33;
  assign _GEN_5749 = {{8'd0}, programBufferMem_33};
  assign _T_5934 = _GEN_5749 << 8;
  assign _GEN_5750 = {{8'd0}, programBufferMem_32};
  assign _T_5938 = _GEN_5750 | _T_5934;
  assign _T_5954 = _T_7458 & _T_3661;
  assign _T_5958 = _T_7755 & _T_3665;
  assign _GEN_116 = _T_5958 ? _T_3679 : programBufferMem_34;
  assign _GEN_5751 = {{16'd0}, programBufferMem_34};
  assign _T_5974 = _GEN_5751 << 16;
  assign _GEN_5752 = {{8'd0}, _T_5938};
  assign _T_5978 = _GEN_5752 | _T_5974;
  assign _T_5994 = _T_7458 & _T_3701;
  assign _T_5998 = _T_7755 & _T_3705;
  assign _GEN_117 = _T_5998 ? _T_3719 : programBufferMem_35;
  assign _GEN_5753 = {{24'd0}, programBufferMem_35};
  assign _T_6014 = _GEN_5753 << 24;
  assign _GEN_5754 = {{8'd0}, _T_5978};
  assign _T_6018 = _GEN_5754 | _T_6014;
  assign _T_6038 = _T_7619 & _T_3745;
  assign _GEN_118 = _T_6038 ? io_dmi_in_0_a_bits_data : 32'h0;
  assign _T_6074 = _T_7426 & _T_3581;
  assign _T_6078 = _T_7723 & _T_3585;
  assign _GEN_119 = _T_6078 ? _T_3599 : programBufferMem_16;
  assign _T_6114 = _T_7426 & _T_3621;
  assign _T_6118 = _T_7723 & _T_3625;
  assign _GEN_120 = _T_6118 ? _T_3639 : programBufferMem_17;
  assign _GEN_5755 = {{8'd0}, programBufferMem_17};
  assign _T_6134 = _GEN_5755 << 8;
  assign _GEN_5756 = {{8'd0}, programBufferMem_16};
  assign _T_6138 = _GEN_5756 | _T_6134;
  assign _T_6154 = _T_7426 & _T_3661;
  assign _T_6158 = _T_7723 & _T_3665;
  assign _GEN_121 = _T_6158 ? _T_3679 : programBufferMem_18;
  assign _GEN_5757 = {{16'd0}, programBufferMem_18};
  assign _T_6174 = _GEN_5757 << 16;
  assign _GEN_5758 = {{8'd0}, _T_6138};
  assign _T_6178 = _GEN_5758 | _T_6174;
  assign _T_6194 = _T_7426 & _T_3701;
  assign _T_6198 = _T_7723 & _T_3705;
  assign _GEN_122 = _T_6198 ? _T_3719 : programBufferMem_19;
  assign _GEN_5759 = {{24'd0}, programBufferMem_19};
  assign _T_6214 = _GEN_5759 << 24;
  assign _GEN_5760 = {{8'd0}, _T_6178};
  assign _T_6218 = _GEN_5760 | _T_6214;
  assign _T_6274 = _T_7298 & _T_3581;
  assign _T_6278 = _T_7595 & _T_3585;
  assign _GEN_123 = _T_6278 ? _T_3599 : abstractDataMem_0;
  assign _T_6314 = _T_7298 & _T_3621;
  assign _T_6318 = _T_7595 & _T_3625;
  assign _GEN_124 = _T_6318 ? _T_3639 : abstractDataMem_1;
  assign _GEN_5761 = {{8'd0}, abstractDataMem_1};
  assign _T_6334 = _GEN_5761 << 8;
  assign _GEN_5762 = {{8'd0}, abstractDataMem_0};
  assign _T_6338 = _GEN_5762 | _T_6334;
  assign _T_6354 = _T_7298 & _T_3661;
  assign _T_6358 = _T_7595 & _T_3665;
  assign _GEN_125 = _T_6358 ? _T_3679 : abstractDataMem_2;
  assign _GEN_5763 = {{16'd0}, abstractDataMem_2};
  assign _T_6374 = _GEN_5763 << 16;
  assign _GEN_5764 = {{8'd0}, _T_6338};
  assign _T_6378 = _GEN_5764 | _T_6374;
  assign _T_6394 = _T_7298 & _T_3701;
  assign _T_6398 = _T_7595 & _T_3705;
  assign _GEN_126 = _T_6398 ? _T_3719 : abstractDataMem_3;
  assign _GEN_5765 = {{24'd0}, abstractDataMem_3};
  assign _T_6414 = _GEN_5765 << 24;
  assign _GEN_5766 = {{8'd0}, _T_6378};
  assign _T_6418 = _GEN_5766 | _T_6414;
  assign _T_6434 = _T_7514 & _T_3581;
  assign _T_6438 = _T_7811 & _T_3585;
  assign _GEN_127 = _T_6438 ? _T_3599 : programBufferMem_60;
  assign _T_6474 = _T_7514 & _T_3621;
  assign _T_6478 = _T_7811 & _T_3625;
  assign _GEN_128 = _T_6478 ? _T_3639 : programBufferMem_61;
  assign _GEN_5767 = {{8'd0}, programBufferMem_61};
  assign _T_6494 = _GEN_5767 << 8;
  assign _GEN_5768 = {{8'd0}, programBufferMem_60};
  assign _T_6498 = _GEN_5768 | _T_6494;
  assign _T_6514 = _T_7514 & _T_3661;
  assign _T_6518 = _T_7811 & _T_3665;
  assign _GEN_129 = _T_6518 ? _T_3679 : programBufferMem_62;
  assign _GEN_5769 = {{16'd0}, programBufferMem_62};
  assign _T_6534 = _GEN_5769 << 16;
  assign _GEN_5770 = {{8'd0}, _T_6498};
  assign _T_6538 = _GEN_5770 | _T_6534;
  assign _T_6554 = _T_7514 & _T_3701;
  assign _T_6558 = _T_7811 & _T_3705;
  assign _GEN_130 = _T_6558 ? _T_3719 : programBufferMem_63;
  assign _GEN_5771 = {{24'd0}, programBufferMem_63};
  assign _T_6574 = _GEN_5771 << 24;
  assign _GEN_5772 = {{8'd0}, _T_6538};
  assign _T_6578 = _GEN_5772 | _T_6574;
  assign _T_6579 = _T_2875[0];
  assign _T_6580 = _T_2875[1];
  assign _T_6581 = _T_2875[2];
  assign _T_6582 = _T_2875[3];
  assign _T_6584 = _T_2875[5];
  assign _T_6586 = {_T_6580,_T_6579};
  assign _T_6587 = {_T_6584,_T_6582};
  assign _T_6588 = {_T_6587,_T_6581};
  assign _T_6589 = {_T_6588,_T_6586};
  assign _T_6602 = 32'h1 << _T_6589;
  assign _T_6607 = _T_6602[4];
  assign _T_6609 = _T_6602[6];
  assign _T_6610 = _T_6602[7];
  assign _T_6611 = _T_6602[8];
  assign _T_6619 = _T_6602[16];
  assign _T_6620 = _T_6602[17];
  assign _T_6621 = _T_6602[18];
  assign _T_6622 = _T_6602[19];
  assign _T_6623 = _T_6602[20];
  assign _T_6624 = _T_6602[21];
  assign _T_6625 = _T_6602[22];
  assign _T_6626 = _T_6602[23];
  assign _T_6627 = _T_6602[24];
  assign _T_6628 = _T_6602[25];
  assign _T_6629 = _T_6602[26];
  assign _T_6630 = _T_6602[27];
  assign _T_6631 = _T_6602[28];
  assign _T_6632 = _T_6602[29];
  assign _T_6633 = _T_6602[30];
  assign _T_6634 = _T_6602[31];
  assign _T_6669 = io_dmi_in_0_a_valid & io_dmi_in_0_d_ready;
  assign _T_6670 = _T_6669 & _T_2874;
  assign _T_6705 = _T_6670 & _T_6607;
  assign _T_6801 = _T_6670 & _T_6619;
  assign _T_6809 = _T_6670 & _T_6620;
  assign _T_6817 = _T_6670 & _T_6621;
  assign _T_6825 = _T_6670 & _T_6622;
  assign _T_6833 = _T_6670 & _T_6623;
  assign _T_6841 = _T_6670 & _T_6624;
  assign _T_6849 = _T_6670 & _T_6625;
  assign _T_6857 = _T_6670 & _T_6626;
  assign _T_6865 = _T_6670 & _T_6627;
  assign _T_6873 = _T_6670 & _T_6628;
  assign _T_6881 = _T_6670 & _T_6629;
  assign _T_6889 = _T_6670 & _T_6630;
  assign _T_6897 = _T_6670 & _T_6631;
  assign _T_6905 = _T_6670 & _T_6632;
  assign _T_6913 = _T_6670 & _T_6633;
  assign _T_6921 = _T_6670 & _T_6634;
  assign _T_6966 = _T_2874 == 1'h0;
  assign _T_6967 = _T_6669 & _T_6966;
  assign _T_7002 = _T_6967 & _T_6607;
  assign _T_7018 = _T_6967 & _T_6609;
  assign _T_7026 = _T_6967 & _T_6610;
  assign _T_7034 = _T_6967 & _T_6611;
  assign _T_7098 = _T_6967 & _T_6619;
  assign _T_7106 = _T_6967 & _T_6620;
  assign _T_7114 = _T_6967 & _T_6621;
  assign _T_7122 = _T_6967 & _T_6622;
  assign _T_7130 = _T_6967 & _T_6623;
  assign _T_7138 = _T_6967 & _T_6624;
  assign _T_7146 = _T_6967 & _T_6625;
  assign _T_7154 = _T_6967 & _T_6626;
  assign _T_7162 = _T_6967 & _T_6627;
  assign _T_7170 = _T_6967 & _T_6628;
  assign _T_7178 = _T_6967 & _T_6629;
  assign _T_7186 = _T_6967 & _T_6630;
  assign _T_7194 = _T_6967 & _T_6631;
  assign _T_7202 = _T_6967 & _T_6632;
  assign _T_7210 = _T_6967 & _T_6633;
  assign _T_7218 = _T_6967 & _T_6634;
  assign _T_7298 = _T_6705 & _T_3163;
  assign _T_7394 = _T_6801 & _T_3028;
  assign _T_7402 = _T_6809 & _T_3010;
  assign _T_7410 = _T_6817 & _T_3037;
  assign _T_7418 = _T_6825 & _T_3100;
  assign _T_7426 = _T_6833 & _T_3145;
  assign _T_7434 = _T_6841 & _T_2983;
  assign _T_7442 = _T_6849 & _T_3001;
  assign _T_7450 = _T_6857 & _T_3091;
  assign _T_7458 = _T_6865 & _T_3127;
  assign _T_7466 = _T_6873 & _T_3019;
  assign _T_7474 = _T_6881 & _T_2965;
  assign _T_7482 = _T_6889 & _T_3118;
  assign _T_7490 = _T_6897 & _T_3082;
  assign _T_7498 = _T_6905 & _T_3046;
  assign _T_7506 = _T_6913 & _T_2992;
  assign _T_7514 = _T_6921 & _T_3172;
  assign _T_7595 = _T_7002 & _T_3163;
  assign _T_7611 = _T_7018 & _T_3073;
  assign _T_7619 = _T_7026 & _T_3136;
  assign _T_7627 = _T_7034 & _T_2974;
  assign _T_7691 = _T_7098 & _T_3028;
  assign _T_7699 = _T_7106 & _T_3010;
  assign _T_7707 = _T_7114 & _T_3037;
  assign _T_7715 = _T_7122 & _T_3100;
  assign _T_7723 = _T_7130 & _T_3145;
  assign _T_7731 = _T_7138 & _T_2983;
  assign _T_7739 = _T_7146 & _T_3001;
  assign _T_7747 = _T_7154 & _T_3091;
  assign _T_7755 = _T_7162 & _T_3127;
  assign _T_7763 = _T_7170 & _T_3019;
  assign _T_7771 = _T_7178 & _T_2965;
  assign _T_7779 = _T_7186 & _T_3118;
  assign _T_7787 = _T_7194 & _T_3082;
  assign _T_7795 = _T_7202 & _T_3046;
  assign _T_7803 = _T_7210 & _T_2992;
  assign _T_7811 = _T_7218 & _T_3172;
  assign _GEN_255 = 5'h1 == _T_6589 ? _T_3064 : _T_3055;
  assign _GEN_256 = 5'h2 == _T_6589 ? _T_3109 : _GEN_255;
  assign _GEN_257 = 5'h3 == _T_6589 ? _T_3154 : _GEN_256;
  assign _GEN_258 = 5'h4 == _T_6589 ? _T_3163 : _GEN_257;
  assign _GEN_259 = 5'h5 == _T_6589 ? 1'h1 : _GEN_258;
  assign _GEN_260 = 5'h6 == _T_6589 ? _T_3073 : _GEN_259;
  assign _GEN_261 = 5'h7 == _T_6589 ? _T_3136 : _GEN_260;
  assign _GEN_262 = 5'h8 == _T_6589 ? _T_2974 : _GEN_261;
  assign _GEN_263 = 5'h9 == _T_6589 ? 1'h1 : _GEN_262;
  assign _GEN_264 = 5'ha == _T_6589 ? 1'h1 : _GEN_263;
  assign _GEN_265 = 5'hb == _T_6589 ? 1'h1 : _GEN_264;
  assign _GEN_266 = 5'hc == _T_6589 ? 1'h1 : _GEN_265;
  assign _GEN_267 = 5'hd == _T_6589 ? 1'h1 : _GEN_266;
  assign _GEN_268 = 5'he == _T_6589 ? 1'h1 : _GEN_267;
  assign _GEN_269 = 5'hf == _T_6589 ? 1'h1 : _GEN_268;
  assign _GEN_270 = 5'h10 == _T_6589 ? _T_3028 : _GEN_269;
  assign _GEN_271 = 5'h11 == _T_6589 ? _T_3010 : _GEN_270;
  assign _GEN_272 = 5'h12 == _T_6589 ? _T_3037 : _GEN_271;
  assign _GEN_273 = 5'h13 == _T_6589 ? _T_3100 : _GEN_272;
  assign _GEN_274 = 5'h14 == _T_6589 ? _T_3145 : _GEN_273;
  assign _GEN_275 = 5'h15 == _T_6589 ? _T_2983 : _GEN_274;
  assign _GEN_276 = 5'h16 == _T_6589 ? _T_3001 : _GEN_275;
  assign _GEN_277 = 5'h17 == _T_6589 ? _T_3091 : _GEN_276;
  assign _GEN_278 = 5'h18 == _T_6589 ? _T_3127 : _GEN_277;
  assign _GEN_279 = 5'h19 == _T_6589 ? _T_3019 : _GEN_278;
  assign _GEN_280 = 5'h1a == _T_6589 ? _T_2965 : _GEN_279;
  assign _GEN_281 = 5'h1b == _T_6589 ? _T_3118 : _GEN_280;
  assign _GEN_282 = 5'h1c == _T_6589 ? _T_3082 : _GEN_281;
  assign _GEN_283 = 5'h1d == _T_6589 ? _T_3046 : _GEN_282;
  assign _GEN_284 = 5'h1e == _T_6589 ? _T_2992 : _GEN_283;
  assign _GEN_285 = 5'h1f == _T_6589 ? _T_3172 : _GEN_284;
  assign _GEN_286 = 5'h1 == _T_6589 ? _T_2817 : haltedStatus_0;
  assign _GEN_287 = 5'h2 == _T_6589 ? 32'h111380 : _GEN_286;
  assign _GEN_288 = 5'h3 == _T_6589 ? _T_2853 : _GEN_287;
  assign _GEN_289 = 5'h4 == _T_6589 ? _T_6418 : _GEN_288;
  assign _GEN_290 = 5'h5 == _T_6589 ? 32'h0 : _GEN_289;
  assign _GEN_291 = 5'h6 == _T_6589 ? _T_2860 : _GEN_290;
  assign _GEN_292 = 5'h7 == _T_6589 ? _T_2863 : _GEN_291;
  assign _GEN_293 = 5'h8 == _T_6589 ? _T_2862 : _GEN_292;
  assign _GEN_294 = 5'h9 == _T_6589 ? 32'h0 : _GEN_293;
  assign _GEN_295 = 5'ha == _T_6589 ? 32'h0 : _GEN_294;
  assign _GEN_296 = 5'hb == _T_6589 ? 32'h0 : _GEN_295;
  assign _GEN_297 = 5'hc == _T_6589 ? 32'h0 : _GEN_296;
  assign _GEN_298 = 5'hd == _T_6589 ? 32'h0 : _GEN_297;
  assign _GEN_299 = 5'he == _T_6589 ? 32'h0 : _GEN_298;
  assign _GEN_300 = 5'hf == _T_6589 ? 32'h0 : _GEN_299;
  assign _GEN_301 = 5'h10 == _T_6589 ? _T_4738 : _GEN_300;
  assign _GEN_302 = 5'h11 == _T_6589 ? _T_4418 : _GEN_301;
  assign _GEN_303 = 5'h12 == _T_6589 ? _T_4898 : _GEN_302;
  assign _GEN_304 = 5'h13 == _T_6589 ? _T_5658 : _GEN_303;
  assign _GEN_305 = 5'h14 == _T_6589 ? _T_6218 : _GEN_304;
  assign _GEN_306 = 5'h15 == _T_6589 ? _T_3938 : _GEN_305;
  assign _GEN_307 = 5'h16 == _T_6589 ? _T_4258 : _GEN_306;
  assign _GEN_308 = 5'h17 == _T_6589 ? _T_5498 : _GEN_307;
  assign _GEN_309 = 5'h18 == _T_6589 ? _T_6018 : _GEN_308;
  assign _GEN_310 = 5'h19 == _T_6589 ? _T_4578 : _GEN_309;
  assign _GEN_311 = 5'h1a == _T_6589 ? _T_3738 : _GEN_310;
  assign _GEN_312 = 5'h1b == _T_6589 ? _T_5858 : _GEN_311;
  assign _GEN_313 = 5'h1c == _T_6589 ? _T_5338 : _GEN_312;
  assign _GEN_314 = 5'h1d == _T_6589 ? _T_5058 : _GEN_313;
  assign _GEN_315 = 5'h1e == _T_6589 ? _T_4098 : _GEN_314;
  assign _GEN_316 = 5'h1f == _T_6589 ? _T_6578 : _GEN_315;
  assign _T_7940 = _GEN_285 ? _GEN_316 : 32'h0;
  assign _T_7941 = _T_2876[2];
  assign _T_7942 = _T_2876[1:0];
  assign _T_7956 = _T_6278 & _T_103519;
  assign _GEN_317 = _T_7956 ? _GEN_123 : abstractDataMem_0;
  assign _T_7957 = _T_6318 & _T_103519;
  assign _GEN_318 = _T_7957 ? _GEN_124 : abstractDataMem_1;
  assign _T_7958 = _T_6358 & _T_103519;
  assign _GEN_319 = _T_7958 ? _GEN_125 : abstractDataMem_2;
  assign _T_7959 = _T_6398 & _T_103519;
  assign _GEN_320 = _T_7959 ? _GEN_126 : abstractDataMem_3;
  assign _T_7960 = _T_4598 & _T_103521;
  assign _GEN_321 = _T_7960 ? _GEN_85 : programBufferMem_0;
  assign _T_7961 = _T_4638 & _T_103521;
  assign _GEN_322 = _T_7961 ? _GEN_86 : programBufferMem_1;
  assign _T_7962 = _T_4678 & _T_103521;
  assign _GEN_323 = _T_7962 ? _GEN_87 : programBufferMem_2;
  assign _T_7963 = _T_4718 & _T_103521;
  assign _GEN_324 = _T_7963 ? _GEN_88 : programBufferMem_3;
  assign _T_7964 = _T_4278 & _T_103521;
  assign _GEN_325 = _T_7964 ? _GEN_77 : programBufferMem_4;
  assign _T_7965 = _T_4318 & _T_103521;
  assign _GEN_326 = _T_7965 ? _GEN_78 : programBufferMem_5;
  assign _T_7966 = _T_4358 & _T_103521;
  assign _GEN_327 = _T_7966 ? _GEN_79 : programBufferMem_6;
  assign _T_7967 = _T_4398 & _T_103521;
  assign _GEN_328 = _T_7967 ? _GEN_80 : programBufferMem_7;
  assign _T_7968 = _T_4758 & _T_103521;
  assign _GEN_329 = _T_7968 ? _GEN_89 : programBufferMem_8;
  assign _T_7969 = _T_4798 & _T_103521;
  assign _GEN_330 = _T_7969 ? _GEN_90 : programBufferMem_9;
  assign _T_7970 = _T_4838 & _T_103521;
  assign _GEN_331 = _T_7970 ? _GEN_91 : programBufferMem_10;
  assign _T_7971 = _T_4878 & _T_103521;
  assign _GEN_332 = _T_7971 ? _GEN_92 : programBufferMem_11;
  assign _T_7972 = _T_5518 & _T_103521;
  assign _GEN_333 = _T_7972 ? _GEN_106 : programBufferMem_12;
  assign _T_7973 = _T_5558 & _T_103521;
  assign _GEN_334 = _T_7973 ? _GEN_107 : programBufferMem_13;
  assign _T_7974 = _T_5598 & _T_103521;
  assign _GEN_335 = _T_7974 ? _GEN_108 : programBufferMem_14;
  assign _T_7975 = _T_5638 & _T_103521;
  assign _GEN_336 = _T_7975 ? _GEN_109 : programBufferMem_15;
  assign _T_7976 = _T_6078 & _T_103521;
  assign _GEN_337 = _T_7976 ? _GEN_119 : programBufferMem_16;
  assign _T_7977 = _T_6118 & _T_103521;
  assign _GEN_338 = _T_7977 ? _GEN_120 : programBufferMem_17;
  assign _T_7978 = _T_6158 & _T_103521;
  assign _GEN_339 = _T_7978 ? _GEN_121 : programBufferMem_18;
  assign _T_7979 = _T_6198 & _T_103521;
  assign _GEN_340 = _T_7979 ? _GEN_122 : programBufferMem_19;
  assign _T_7980 = _T_3798 & _T_103521;
  assign _GEN_341 = _T_7980 ? _GEN_65 : programBufferMem_20;
  assign _T_7981 = _T_3838 & _T_103521;
  assign _GEN_342 = _T_7981 ? _GEN_66 : programBufferMem_21;
  assign _T_7982 = _T_3878 & _T_103521;
  assign _GEN_343 = _T_7982 ? _GEN_67 : programBufferMem_22;
  assign _T_7983 = _T_3918 & _T_103521;
  assign _GEN_344 = _T_7983 ? _GEN_68 : programBufferMem_23;
  assign _T_7984 = _T_4118 & _T_103521;
  assign _GEN_345 = _T_7984 ? _GEN_73 : programBufferMem_24;
  assign _T_7985 = _T_4158 & _T_103521;
  assign _GEN_346 = _T_7985 ? _GEN_74 : programBufferMem_25;
  assign _T_7986 = _T_4198 & _T_103521;
  assign _GEN_347 = _T_7986 ? _GEN_75 : programBufferMem_26;
  assign _T_7987 = _T_4238 & _T_103521;
  assign _GEN_348 = _T_7987 ? _GEN_76 : programBufferMem_27;
  assign _T_7988 = _T_5358 & _T_103521;
  assign _GEN_349 = _T_7988 ? _GEN_102 : programBufferMem_28;
  assign _T_7989 = _T_5398 & _T_103521;
  assign _GEN_350 = _T_7989 ? _GEN_103 : programBufferMem_29;
  assign _T_7990 = _T_5438 & _T_103521;
  assign _GEN_351 = _T_7990 ? _GEN_104 : programBufferMem_30;
  assign _T_7991 = _T_5478 & _T_103521;
  assign _GEN_352 = _T_7991 ? _GEN_105 : programBufferMem_31;
  assign _T_7992 = _T_5878 & _T_103521;
  assign _GEN_353 = _T_7992 ? _GEN_114 : programBufferMem_32;
  assign _T_7993 = _T_5918 & _T_103521;
  assign _GEN_354 = _T_7993 ? _GEN_115 : programBufferMem_33;
  assign _T_7994 = _T_5958 & _T_103521;
  assign _GEN_355 = _T_7994 ? _GEN_116 : programBufferMem_34;
  assign _T_7995 = _T_5998 & _T_103521;
  assign _GEN_356 = _T_7995 ? _GEN_117 : programBufferMem_35;
  assign _T_7996 = _T_4438 & _T_103521;
  assign _GEN_357 = _T_7996 ? _GEN_81 : programBufferMem_36;
  assign _T_7997 = _T_4478 & _T_103521;
  assign _GEN_358 = _T_7997 ? _GEN_82 : programBufferMem_37;
  assign _T_7998 = _T_4518 & _T_103521;
  assign _GEN_359 = _T_7998 ? _GEN_83 : programBufferMem_38;
  assign _T_7999 = _T_4558 & _T_103521;
  assign _GEN_360 = _T_7999 ? _GEN_84 : programBufferMem_39;
  assign _T_8000 = _T_3598 & _T_103521;
  assign _GEN_361 = _T_8000 ? _GEN_60 : programBufferMem_40;
  assign _T_8001 = _T_3638 & _T_103521;
  assign _GEN_362 = _T_8001 ? _GEN_61 : programBufferMem_41;
  assign _T_8002 = _T_3678 & _T_103521;
  assign _GEN_363 = _T_8002 ? _GEN_62 : programBufferMem_42;
  assign _T_8003 = _T_3718 & _T_103521;
  assign _GEN_364 = _T_8003 ? _GEN_63 : programBufferMem_43;
  assign _T_8004 = _T_5718 & _T_103521;
  assign _GEN_365 = _T_8004 ? _GEN_110 : programBufferMem_44;
  assign _T_8005 = _T_5758 & _T_103521;
  assign _GEN_366 = _T_8005 ? _GEN_111 : programBufferMem_45;
  assign _T_8006 = _T_5798 & _T_103521;
  assign _GEN_367 = _T_8006 ? _GEN_112 : programBufferMem_46;
  assign _T_8007 = _T_5838 & _T_103521;
  assign _GEN_368 = _T_8007 ? _GEN_113 : programBufferMem_47;
  assign _T_8008 = _T_5198 & _T_103521;
  assign _GEN_369 = _T_8008 ? _GEN_98 : programBufferMem_48;
  assign _T_8009 = _T_5238 & _T_103521;
  assign _GEN_370 = _T_8009 ? _GEN_99 : programBufferMem_49;
  assign _T_8010 = _T_5278 & _T_103521;
  assign _GEN_371 = _T_8010 ? _GEN_100 : programBufferMem_50;
  assign _T_8011 = _T_5318 & _T_103521;
  assign _GEN_372 = _T_8011 ? _GEN_101 : programBufferMem_51;
  assign _T_8012 = _T_4918 & _T_103521;
  assign _GEN_373 = _T_8012 ? _GEN_93 : programBufferMem_52;
  assign _T_8013 = _T_4958 & _T_103521;
  assign _GEN_374 = _T_8013 ? _GEN_94 : programBufferMem_53;
  assign _T_8014 = _T_4998 & _T_103521;
  assign _GEN_375 = _T_8014 ? _GEN_95 : programBufferMem_54;
  assign _T_8015 = _T_5038 & _T_103521;
  assign _GEN_376 = _T_8015 ? _GEN_96 : programBufferMem_55;
  assign _T_8016 = _T_3958 & _T_103521;
  assign _GEN_377 = _T_8016 ? _GEN_69 : programBufferMem_56;
  assign _T_8017 = _T_3998 & _T_103521;
  assign _GEN_378 = _T_8017 ? _GEN_70 : programBufferMem_57;
  assign _T_8018 = _T_4038 & _T_103521;
  assign _GEN_379 = _T_8018 ? _GEN_71 : programBufferMem_58;
  assign _T_8019 = _T_4078 & _T_103521;
  assign _GEN_380 = _T_8019 ? _GEN_72 : programBufferMem_59;
  assign _T_8020 = _T_6438 & _T_103521;
  assign _GEN_381 = _T_8020 ? _GEN_127 : programBufferMem_60;
  assign _T_8021 = _T_6478 & _T_103521;
  assign _GEN_382 = _T_8021 ? _GEN_128 : programBufferMem_61;
  assign _T_8022 = _T_6518 & _T_103521;
  assign _GEN_383 = _T_8022 ? _GEN_129 : programBufferMem_62;
  assign _T_8023 = _T_6558 & _T_103521;
  assign _GEN_384 = _T_8023 ? _GEN_130 : programBufferMem_63;
  assign _GEN_385 = _T_1403 ? 1'h0 : goReg;
  assign _GEN_386 = _GEN_5663 ? 1'h1 : _GEN_385;
  assign _T_8235 = _GEN_5663 == 1'h0;
  assign _T_8236 = _T_8235 & _T_50183;
  assign _T_8238 = _T_50184 == 10'h0;
  assign _T_8239 = _T_8238 | reset;
  assign _T_8241 = _T_8239 == 1'h0;
  assign _GEN_387 = _T_8236 ? 1'h0 : _GEN_386;
  assign _GEN_388 = _T_1405 ? _GEN_387 : _GEN_385;
  assign _GEN_389 = 10'h0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_390 = 10'h1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_391 = 10'h2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_392 = 10'h3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_393 = 10'h4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_394 = 10'h5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_395 = 10'h6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_396 = 10'h7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_397 = 10'h8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_398 = 10'h9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_399 = 10'ha == selectedHartReg ? goReg : 1'h0;
  assign _GEN_400 = 10'hb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_401 = 10'hc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_402 = 10'hd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_403 = 10'he == selectedHartReg ? goReg : 1'h0;
  assign _GEN_404 = 10'hf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_405 = 10'h10 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_406 = 10'h11 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_407 = 10'h12 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_408 = 10'h13 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_409 = 10'h14 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_410 = 10'h15 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_411 = 10'h16 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_412 = 10'h17 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_413 = 10'h18 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_414 = 10'h19 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_415 = 10'h1a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_416 = 10'h1b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_417 = 10'h1c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_418 = 10'h1d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_419 = 10'h1e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_420 = 10'h1f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_421 = 10'h20 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_422 = 10'h21 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_423 = 10'h22 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_424 = 10'h23 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_425 = 10'h24 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_426 = 10'h25 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_427 = 10'h26 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_428 = 10'h27 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_429 = 10'h28 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_430 = 10'h29 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_431 = 10'h2a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_432 = 10'h2b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_433 = 10'h2c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_434 = 10'h2d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_435 = 10'h2e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_436 = 10'h2f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_437 = 10'h30 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_438 = 10'h31 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_439 = 10'h32 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_440 = 10'h33 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_441 = 10'h34 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_442 = 10'h35 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_443 = 10'h36 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_444 = 10'h37 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_445 = 10'h38 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_446 = 10'h39 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_447 = 10'h3a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_448 = 10'h3b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_449 = 10'h3c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_450 = 10'h3d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_451 = 10'h3e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_452 = 10'h3f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_453 = 10'h40 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_454 = 10'h41 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_455 = 10'h42 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_456 = 10'h43 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_457 = 10'h44 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_458 = 10'h45 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_459 = 10'h46 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_460 = 10'h47 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_461 = 10'h48 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_462 = 10'h49 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_463 = 10'h4a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_464 = 10'h4b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_465 = 10'h4c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_466 = 10'h4d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_467 = 10'h4e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_468 = 10'h4f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_469 = 10'h50 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_470 = 10'h51 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_471 = 10'h52 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_472 = 10'h53 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_473 = 10'h54 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_474 = 10'h55 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_475 = 10'h56 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_476 = 10'h57 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_477 = 10'h58 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_478 = 10'h59 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_479 = 10'h5a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_480 = 10'h5b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_481 = 10'h5c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_482 = 10'h5d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_483 = 10'h5e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_484 = 10'h5f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_485 = 10'h60 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_486 = 10'h61 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_487 = 10'h62 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_488 = 10'h63 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_489 = 10'h64 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_490 = 10'h65 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_491 = 10'h66 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_492 = 10'h67 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_493 = 10'h68 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_494 = 10'h69 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_495 = 10'h6a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_496 = 10'h6b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_497 = 10'h6c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_498 = 10'h6d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_499 = 10'h6e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_500 = 10'h6f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_501 = 10'h70 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_502 = 10'h71 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_503 = 10'h72 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_504 = 10'h73 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_505 = 10'h74 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_506 = 10'h75 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_507 = 10'h76 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_508 = 10'h77 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_509 = 10'h78 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_510 = 10'h79 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_511 = 10'h7a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_512 = 10'h7b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_513 = 10'h7c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_514 = 10'h7d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_515 = 10'h7e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_516 = 10'h7f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_517 = 10'h80 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_518 = 10'h81 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_519 = 10'h82 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_520 = 10'h83 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_521 = 10'h84 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_522 = 10'h85 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_523 = 10'h86 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_524 = 10'h87 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_525 = 10'h88 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_526 = 10'h89 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_527 = 10'h8a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_528 = 10'h8b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_529 = 10'h8c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_530 = 10'h8d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_531 = 10'h8e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_532 = 10'h8f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_533 = 10'h90 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_534 = 10'h91 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_535 = 10'h92 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_536 = 10'h93 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_537 = 10'h94 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_538 = 10'h95 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_539 = 10'h96 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_540 = 10'h97 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_541 = 10'h98 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_542 = 10'h99 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_543 = 10'h9a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_544 = 10'h9b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_545 = 10'h9c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_546 = 10'h9d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_547 = 10'h9e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_548 = 10'h9f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_549 = 10'ha0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_550 = 10'ha1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_551 = 10'ha2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_552 = 10'ha3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_553 = 10'ha4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_554 = 10'ha5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_555 = 10'ha6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_556 = 10'ha7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_557 = 10'ha8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_558 = 10'ha9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_559 = 10'haa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_560 = 10'hab == selectedHartReg ? goReg : 1'h0;
  assign _GEN_561 = 10'hac == selectedHartReg ? goReg : 1'h0;
  assign _GEN_562 = 10'had == selectedHartReg ? goReg : 1'h0;
  assign _GEN_563 = 10'hae == selectedHartReg ? goReg : 1'h0;
  assign _GEN_564 = 10'haf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_565 = 10'hb0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_566 = 10'hb1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_567 = 10'hb2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_568 = 10'hb3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_569 = 10'hb4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_570 = 10'hb5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_571 = 10'hb6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_572 = 10'hb7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_573 = 10'hb8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_574 = 10'hb9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_575 = 10'hba == selectedHartReg ? goReg : 1'h0;
  assign _GEN_576 = 10'hbb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_577 = 10'hbc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_578 = 10'hbd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_579 = 10'hbe == selectedHartReg ? goReg : 1'h0;
  assign _GEN_580 = 10'hbf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_581 = 10'hc0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_582 = 10'hc1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_583 = 10'hc2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_584 = 10'hc3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_585 = 10'hc4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_586 = 10'hc5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_587 = 10'hc6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_588 = 10'hc7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_589 = 10'hc8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_590 = 10'hc9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_591 = 10'hca == selectedHartReg ? goReg : 1'h0;
  assign _GEN_592 = 10'hcb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_593 = 10'hcc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_594 = 10'hcd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_595 = 10'hce == selectedHartReg ? goReg : 1'h0;
  assign _GEN_596 = 10'hcf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_597 = 10'hd0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_598 = 10'hd1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_599 = 10'hd2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_600 = 10'hd3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_601 = 10'hd4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_602 = 10'hd5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_603 = 10'hd6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_604 = 10'hd7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_605 = 10'hd8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_606 = 10'hd9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_607 = 10'hda == selectedHartReg ? goReg : 1'h0;
  assign _GEN_608 = 10'hdb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_609 = 10'hdc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_610 = 10'hdd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_611 = 10'hde == selectedHartReg ? goReg : 1'h0;
  assign _GEN_612 = 10'hdf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_613 = 10'he0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_614 = 10'he1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_615 = 10'he2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_616 = 10'he3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_617 = 10'he4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_618 = 10'he5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_619 = 10'he6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_620 = 10'he7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_621 = 10'he8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_622 = 10'he9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_623 = 10'hea == selectedHartReg ? goReg : 1'h0;
  assign _GEN_624 = 10'heb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_625 = 10'hec == selectedHartReg ? goReg : 1'h0;
  assign _GEN_626 = 10'hed == selectedHartReg ? goReg : 1'h0;
  assign _GEN_627 = 10'hee == selectedHartReg ? goReg : 1'h0;
  assign _GEN_628 = 10'hef == selectedHartReg ? goReg : 1'h0;
  assign _GEN_629 = 10'hf0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_630 = 10'hf1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_631 = 10'hf2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_632 = 10'hf3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_633 = 10'hf4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_634 = 10'hf5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_635 = 10'hf6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_636 = 10'hf7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_637 = 10'hf8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_638 = 10'hf9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_639 = 10'hfa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_640 = 10'hfb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_641 = 10'hfc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_642 = 10'hfd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_643 = 10'hfe == selectedHartReg ? goReg : 1'h0;
  assign _GEN_644 = 10'hff == selectedHartReg ? goReg : 1'h0;
  assign _GEN_645 = 10'h100 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_646 = 10'h101 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_647 = 10'h102 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_648 = 10'h103 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_649 = 10'h104 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_650 = 10'h105 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_651 = 10'h106 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_652 = 10'h107 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_653 = 10'h108 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_654 = 10'h109 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_655 = 10'h10a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_656 = 10'h10b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_657 = 10'h10c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_658 = 10'h10d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_659 = 10'h10e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_660 = 10'h10f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_661 = 10'h110 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_662 = 10'h111 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_663 = 10'h112 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_664 = 10'h113 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_665 = 10'h114 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_666 = 10'h115 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_667 = 10'h116 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_668 = 10'h117 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_669 = 10'h118 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_670 = 10'h119 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_671 = 10'h11a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_672 = 10'h11b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_673 = 10'h11c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_674 = 10'h11d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_675 = 10'h11e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_676 = 10'h11f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_677 = 10'h120 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_678 = 10'h121 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_679 = 10'h122 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_680 = 10'h123 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_681 = 10'h124 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_682 = 10'h125 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_683 = 10'h126 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_684 = 10'h127 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_685 = 10'h128 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_686 = 10'h129 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_687 = 10'h12a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_688 = 10'h12b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_689 = 10'h12c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_690 = 10'h12d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_691 = 10'h12e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_692 = 10'h12f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_693 = 10'h130 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_694 = 10'h131 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_695 = 10'h132 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_696 = 10'h133 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_697 = 10'h134 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_698 = 10'h135 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_699 = 10'h136 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_700 = 10'h137 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_701 = 10'h138 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_702 = 10'h139 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_703 = 10'h13a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_704 = 10'h13b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_705 = 10'h13c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_706 = 10'h13d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_707 = 10'h13e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_708 = 10'h13f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_709 = 10'h140 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_710 = 10'h141 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_711 = 10'h142 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_712 = 10'h143 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_713 = 10'h144 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_714 = 10'h145 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_715 = 10'h146 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_716 = 10'h147 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_717 = 10'h148 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_718 = 10'h149 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_719 = 10'h14a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_720 = 10'h14b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_721 = 10'h14c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_722 = 10'h14d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_723 = 10'h14e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_724 = 10'h14f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_725 = 10'h150 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_726 = 10'h151 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_727 = 10'h152 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_728 = 10'h153 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_729 = 10'h154 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_730 = 10'h155 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_731 = 10'h156 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_732 = 10'h157 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_733 = 10'h158 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_734 = 10'h159 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_735 = 10'h15a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_736 = 10'h15b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_737 = 10'h15c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_738 = 10'h15d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_739 = 10'h15e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_740 = 10'h15f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_741 = 10'h160 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_742 = 10'h161 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_743 = 10'h162 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_744 = 10'h163 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_745 = 10'h164 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_746 = 10'h165 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_747 = 10'h166 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_748 = 10'h167 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_749 = 10'h168 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_750 = 10'h169 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_751 = 10'h16a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_752 = 10'h16b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_753 = 10'h16c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_754 = 10'h16d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_755 = 10'h16e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_756 = 10'h16f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_757 = 10'h170 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_758 = 10'h171 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_759 = 10'h172 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_760 = 10'h173 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_761 = 10'h174 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_762 = 10'h175 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_763 = 10'h176 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_764 = 10'h177 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_765 = 10'h178 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_766 = 10'h179 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_767 = 10'h17a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_768 = 10'h17b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_769 = 10'h17c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_770 = 10'h17d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_771 = 10'h17e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_772 = 10'h17f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_773 = 10'h180 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_774 = 10'h181 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_775 = 10'h182 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_776 = 10'h183 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_777 = 10'h184 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_778 = 10'h185 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_779 = 10'h186 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_780 = 10'h187 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_781 = 10'h188 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_782 = 10'h189 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_783 = 10'h18a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_784 = 10'h18b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_785 = 10'h18c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_786 = 10'h18d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_787 = 10'h18e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_788 = 10'h18f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_789 = 10'h190 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_790 = 10'h191 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_791 = 10'h192 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_792 = 10'h193 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_793 = 10'h194 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_794 = 10'h195 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_795 = 10'h196 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_796 = 10'h197 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_797 = 10'h198 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_798 = 10'h199 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_799 = 10'h19a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_800 = 10'h19b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_801 = 10'h19c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_802 = 10'h19d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_803 = 10'h19e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_804 = 10'h19f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_805 = 10'h1a0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_806 = 10'h1a1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_807 = 10'h1a2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_808 = 10'h1a3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_809 = 10'h1a4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_810 = 10'h1a5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_811 = 10'h1a6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_812 = 10'h1a7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_813 = 10'h1a8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_814 = 10'h1a9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_815 = 10'h1aa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_816 = 10'h1ab == selectedHartReg ? goReg : 1'h0;
  assign _GEN_817 = 10'h1ac == selectedHartReg ? goReg : 1'h0;
  assign _GEN_818 = 10'h1ad == selectedHartReg ? goReg : 1'h0;
  assign _GEN_819 = 10'h1ae == selectedHartReg ? goReg : 1'h0;
  assign _GEN_820 = 10'h1af == selectedHartReg ? goReg : 1'h0;
  assign _GEN_821 = 10'h1b0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_822 = 10'h1b1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_823 = 10'h1b2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_824 = 10'h1b3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_825 = 10'h1b4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_826 = 10'h1b5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_827 = 10'h1b6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_828 = 10'h1b7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_829 = 10'h1b8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_830 = 10'h1b9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_831 = 10'h1ba == selectedHartReg ? goReg : 1'h0;
  assign _GEN_832 = 10'h1bb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_833 = 10'h1bc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_834 = 10'h1bd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_835 = 10'h1be == selectedHartReg ? goReg : 1'h0;
  assign _GEN_836 = 10'h1bf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_837 = 10'h1c0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_838 = 10'h1c1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_839 = 10'h1c2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_840 = 10'h1c3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_841 = 10'h1c4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_842 = 10'h1c5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_843 = 10'h1c6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_844 = 10'h1c7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_845 = 10'h1c8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_846 = 10'h1c9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_847 = 10'h1ca == selectedHartReg ? goReg : 1'h0;
  assign _GEN_848 = 10'h1cb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_849 = 10'h1cc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_850 = 10'h1cd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_851 = 10'h1ce == selectedHartReg ? goReg : 1'h0;
  assign _GEN_852 = 10'h1cf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_853 = 10'h1d0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_854 = 10'h1d1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_855 = 10'h1d2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_856 = 10'h1d3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_857 = 10'h1d4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_858 = 10'h1d5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_859 = 10'h1d6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_860 = 10'h1d7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_861 = 10'h1d8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_862 = 10'h1d9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_863 = 10'h1da == selectedHartReg ? goReg : 1'h0;
  assign _GEN_864 = 10'h1db == selectedHartReg ? goReg : 1'h0;
  assign _GEN_865 = 10'h1dc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_866 = 10'h1dd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_867 = 10'h1de == selectedHartReg ? goReg : 1'h0;
  assign _GEN_868 = 10'h1df == selectedHartReg ? goReg : 1'h0;
  assign _GEN_869 = 10'h1e0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_870 = 10'h1e1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_871 = 10'h1e2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_872 = 10'h1e3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_873 = 10'h1e4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_874 = 10'h1e5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_875 = 10'h1e6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_876 = 10'h1e7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_877 = 10'h1e8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_878 = 10'h1e9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_879 = 10'h1ea == selectedHartReg ? goReg : 1'h0;
  assign _GEN_880 = 10'h1eb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_881 = 10'h1ec == selectedHartReg ? goReg : 1'h0;
  assign _GEN_882 = 10'h1ed == selectedHartReg ? goReg : 1'h0;
  assign _GEN_883 = 10'h1ee == selectedHartReg ? goReg : 1'h0;
  assign _GEN_884 = 10'h1ef == selectedHartReg ? goReg : 1'h0;
  assign _GEN_885 = 10'h1f0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_886 = 10'h1f1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_887 = 10'h1f2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_888 = 10'h1f3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_889 = 10'h1f4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_890 = 10'h1f5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_891 = 10'h1f6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_892 = 10'h1f7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_893 = 10'h1f8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_894 = 10'h1f9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_895 = 10'h1fa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_896 = 10'h1fb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_897 = 10'h1fc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_898 = 10'h1fd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_899 = 10'h1fe == selectedHartReg ? goReg : 1'h0;
  assign _GEN_900 = 10'h1ff == selectedHartReg ? goReg : 1'h0;
  assign _GEN_901 = 10'h200 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_902 = 10'h201 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_903 = 10'h202 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_904 = 10'h203 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_905 = 10'h204 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_906 = 10'h205 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_907 = 10'h206 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_908 = 10'h207 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_909 = 10'h208 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_910 = 10'h209 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_911 = 10'h20a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_912 = 10'h20b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_913 = 10'h20c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_914 = 10'h20d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_915 = 10'h20e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_916 = 10'h20f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_917 = 10'h210 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_918 = 10'h211 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_919 = 10'h212 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_920 = 10'h213 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_921 = 10'h214 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_922 = 10'h215 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_923 = 10'h216 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_924 = 10'h217 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_925 = 10'h218 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_926 = 10'h219 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_927 = 10'h21a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_928 = 10'h21b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_929 = 10'h21c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_930 = 10'h21d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_931 = 10'h21e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_932 = 10'h21f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_933 = 10'h220 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_934 = 10'h221 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_935 = 10'h222 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_936 = 10'h223 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_937 = 10'h224 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_938 = 10'h225 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_939 = 10'h226 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_940 = 10'h227 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_941 = 10'h228 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_942 = 10'h229 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_943 = 10'h22a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_944 = 10'h22b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_945 = 10'h22c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_946 = 10'h22d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_947 = 10'h22e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_948 = 10'h22f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_949 = 10'h230 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_950 = 10'h231 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_951 = 10'h232 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_952 = 10'h233 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_953 = 10'h234 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_954 = 10'h235 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_955 = 10'h236 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_956 = 10'h237 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_957 = 10'h238 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_958 = 10'h239 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_959 = 10'h23a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_960 = 10'h23b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_961 = 10'h23c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_962 = 10'h23d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_963 = 10'h23e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_964 = 10'h23f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_965 = 10'h240 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_966 = 10'h241 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_967 = 10'h242 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_968 = 10'h243 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_969 = 10'h244 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_970 = 10'h245 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_971 = 10'h246 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_972 = 10'h247 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_973 = 10'h248 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_974 = 10'h249 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_975 = 10'h24a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_976 = 10'h24b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_977 = 10'h24c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_978 = 10'h24d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_979 = 10'h24e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_980 = 10'h24f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_981 = 10'h250 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_982 = 10'h251 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_983 = 10'h252 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_984 = 10'h253 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_985 = 10'h254 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_986 = 10'h255 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_987 = 10'h256 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_988 = 10'h257 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_989 = 10'h258 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_990 = 10'h259 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_991 = 10'h25a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_992 = 10'h25b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_993 = 10'h25c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_994 = 10'h25d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_995 = 10'h25e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_996 = 10'h25f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_997 = 10'h260 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_998 = 10'h261 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_999 = 10'h262 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1000 = 10'h263 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1001 = 10'h264 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1002 = 10'h265 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1003 = 10'h266 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1004 = 10'h267 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1005 = 10'h268 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1006 = 10'h269 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1007 = 10'h26a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1008 = 10'h26b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1009 = 10'h26c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1010 = 10'h26d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1011 = 10'h26e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1012 = 10'h26f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1013 = 10'h270 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1014 = 10'h271 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1015 = 10'h272 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1016 = 10'h273 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1017 = 10'h274 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1018 = 10'h275 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1019 = 10'h276 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1020 = 10'h277 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1021 = 10'h278 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1022 = 10'h279 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1023 = 10'h27a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1024 = 10'h27b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1025 = 10'h27c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1026 = 10'h27d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1027 = 10'h27e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1028 = 10'h27f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1029 = 10'h280 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1030 = 10'h281 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1031 = 10'h282 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1032 = 10'h283 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1033 = 10'h284 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1034 = 10'h285 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1035 = 10'h286 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1036 = 10'h287 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1037 = 10'h288 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1038 = 10'h289 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1039 = 10'h28a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1040 = 10'h28b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1041 = 10'h28c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1042 = 10'h28d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1043 = 10'h28e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1044 = 10'h28f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1045 = 10'h290 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1046 = 10'h291 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1047 = 10'h292 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1048 = 10'h293 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1049 = 10'h294 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1050 = 10'h295 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1051 = 10'h296 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1052 = 10'h297 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1053 = 10'h298 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1054 = 10'h299 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1055 = 10'h29a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1056 = 10'h29b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1057 = 10'h29c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1058 = 10'h29d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1059 = 10'h29e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1060 = 10'h29f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1061 = 10'h2a0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1062 = 10'h2a1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1063 = 10'h2a2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1064 = 10'h2a3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1065 = 10'h2a4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1066 = 10'h2a5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1067 = 10'h2a6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1068 = 10'h2a7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1069 = 10'h2a8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1070 = 10'h2a9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1071 = 10'h2aa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1072 = 10'h2ab == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1073 = 10'h2ac == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1074 = 10'h2ad == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1075 = 10'h2ae == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1076 = 10'h2af == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1077 = 10'h2b0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1078 = 10'h2b1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1079 = 10'h2b2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1080 = 10'h2b3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1081 = 10'h2b4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1082 = 10'h2b5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1083 = 10'h2b6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1084 = 10'h2b7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1085 = 10'h2b8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1086 = 10'h2b9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1087 = 10'h2ba == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1088 = 10'h2bb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1089 = 10'h2bc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1090 = 10'h2bd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1091 = 10'h2be == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1092 = 10'h2bf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1093 = 10'h2c0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1094 = 10'h2c1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1095 = 10'h2c2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1096 = 10'h2c3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1097 = 10'h2c4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1098 = 10'h2c5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1099 = 10'h2c6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1100 = 10'h2c7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1101 = 10'h2c8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1102 = 10'h2c9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1103 = 10'h2ca == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1104 = 10'h2cb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1105 = 10'h2cc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1106 = 10'h2cd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1107 = 10'h2ce == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1108 = 10'h2cf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1109 = 10'h2d0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1110 = 10'h2d1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1111 = 10'h2d2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1112 = 10'h2d3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1113 = 10'h2d4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1114 = 10'h2d5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1115 = 10'h2d6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1116 = 10'h2d7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1117 = 10'h2d8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1118 = 10'h2d9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1119 = 10'h2da == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1120 = 10'h2db == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1121 = 10'h2dc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1122 = 10'h2dd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1123 = 10'h2de == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1124 = 10'h2df == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1125 = 10'h2e0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1126 = 10'h2e1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1127 = 10'h2e2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1128 = 10'h2e3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1129 = 10'h2e4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1130 = 10'h2e5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1131 = 10'h2e6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1132 = 10'h2e7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1133 = 10'h2e8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1134 = 10'h2e9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1135 = 10'h2ea == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1136 = 10'h2eb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1137 = 10'h2ec == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1138 = 10'h2ed == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1139 = 10'h2ee == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1140 = 10'h2ef == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1141 = 10'h2f0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1142 = 10'h2f1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1143 = 10'h2f2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1144 = 10'h2f3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1145 = 10'h2f4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1146 = 10'h2f5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1147 = 10'h2f6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1148 = 10'h2f7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1149 = 10'h2f8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1150 = 10'h2f9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1151 = 10'h2fa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1152 = 10'h2fb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1153 = 10'h2fc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1154 = 10'h2fd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1155 = 10'h2fe == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1156 = 10'h2ff == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1157 = 10'h300 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1158 = 10'h301 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1159 = 10'h302 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1160 = 10'h303 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1161 = 10'h304 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1162 = 10'h305 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1163 = 10'h306 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1164 = 10'h307 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1165 = 10'h308 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1166 = 10'h309 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1167 = 10'h30a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1168 = 10'h30b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1169 = 10'h30c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1170 = 10'h30d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1171 = 10'h30e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1172 = 10'h30f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1173 = 10'h310 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1174 = 10'h311 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1175 = 10'h312 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1176 = 10'h313 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1177 = 10'h314 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1178 = 10'h315 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1179 = 10'h316 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1180 = 10'h317 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1181 = 10'h318 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1182 = 10'h319 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1183 = 10'h31a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1184 = 10'h31b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1185 = 10'h31c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1186 = 10'h31d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1187 = 10'h31e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1188 = 10'h31f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1189 = 10'h320 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1190 = 10'h321 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1191 = 10'h322 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1192 = 10'h323 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1193 = 10'h324 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1194 = 10'h325 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1195 = 10'h326 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1196 = 10'h327 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1197 = 10'h328 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1198 = 10'h329 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1199 = 10'h32a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1200 = 10'h32b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1201 = 10'h32c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1202 = 10'h32d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1203 = 10'h32e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1204 = 10'h32f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1205 = 10'h330 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1206 = 10'h331 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1207 = 10'h332 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1208 = 10'h333 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1209 = 10'h334 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1210 = 10'h335 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1211 = 10'h336 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1212 = 10'h337 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1213 = 10'h338 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1214 = 10'h339 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1215 = 10'h33a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1216 = 10'h33b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1217 = 10'h33c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1218 = 10'h33d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1219 = 10'h33e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1220 = 10'h33f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1221 = 10'h340 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1222 = 10'h341 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1223 = 10'h342 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1224 = 10'h343 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1225 = 10'h344 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1226 = 10'h345 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1227 = 10'h346 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1228 = 10'h347 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1229 = 10'h348 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1230 = 10'h349 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1231 = 10'h34a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1232 = 10'h34b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1233 = 10'h34c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1234 = 10'h34d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1235 = 10'h34e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1236 = 10'h34f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1237 = 10'h350 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1238 = 10'h351 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1239 = 10'h352 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1240 = 10'h353 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1241 = 10'h354 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1242 = 10'h355 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1243 = 10'h356 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1244 = 10'h357 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1245 = 10'h358 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1246 = 10'h359 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1247 = 10'h35a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1248 = 10'h35b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1249 = 10'h35c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1250 = 10'h35d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1251 = 10'h35e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1252 = 10'h35f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1253 = 10'h360 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1254 = 10'h361 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1255 = 10'h362 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1256 = 10'h363 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1257 = 10'h364 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1258 = 10'h365 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1259 = 10'h366 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1260 = 10'h367 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1261 = 10'h368 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1262 = 10'h369 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1263 = 10'h36a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1264 = 10'h36b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1265 = 10'h36c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1266 = 10'h36d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1267 = 10'h36e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1268 = 10'h36f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1269 = 10'h370 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1270 = 10'h371 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1271 = 10'h372 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1272 = 10'h373 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1273 = 10'h374 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1274 = 10'h375 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1275 = 10'h376 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1276 = 10'h377 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1277 = 10'h378 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1278 = 10'h379 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1279 = 10'h37a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1280 = 10'h37b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1281 = 10'h37c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1282 = 10'h37d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1283 = 10'h37e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1284 = 10'h37f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1285 = 10'h380 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1286 = 10'h381 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1287 = 10'h382 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1288 = 10'h383 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1289 = 10'h384 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1290 = 10'h385 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1291 = 10'h386 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1292 = 10'h387 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1293 = 10'h388 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1294 = 10'h389 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1295 = 10'h38a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1296 = 10'h38b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1297 = 10'h38c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1298 = 10'h38d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1299 = 10'h38e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1300 = 10'h38f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1301 = 10'h390 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1302 = 10'h391 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1303 = 10'h392 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1304 = 10'h393 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1305 = 10'h394 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1306 = 10'h395 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1307 = 10'h396 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1308 = 10'h397 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1309 = 10'h398 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1310 = 10'h399 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1311 = 10'h39a == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1312 = 10'h39b == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1313 = 10'h39c == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1314 = 10'h39d == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1315 = 10'h39e == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1316 = 10'h39f == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1317 = 10'h3a0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1318 = 10'h3a1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1319 = 10'h3a2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1320 = 10'h3a3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1321 = 10'h3a4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1322 = 10'h3a5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1323 = 10'h3a6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1324 = 10'h3a7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1325 = 10'h3a8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1326 = 10'h3a9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1327 = 10'h3aa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1328 = 10'h3ab == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1329 = 10'h3ac == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1330 = 10'h3ad == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1331 = 10'h3ae == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1332 = 10'h3af == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1333 = 10'h3b0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1334 = 10'h3b1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1335 = 10'h3b2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1336 = 10'h3b3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1337 = 10'h3b4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1338 = 10'h3b5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1339 = 10'h3b6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1340 = 10'h3b7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1341 = 10'h3b8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1342 = 10'h3b9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1343 = 10'h3ba == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1344 = 10'h3bb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1345 = 10'h3bc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1346 = 10'h3bd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1347 = 10'h3be == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1348 = 10'h3bf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1349 = 10'h3c0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1350 = 10'h3c1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1351 = 10'h3c2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1352 = 10'h3c3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1353 = 10'h3c4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1354 = 10'h3c5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1355 = 10'h3c6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1356 = 10'h3c7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1357 = 10'h3c8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1358 = 10'h3c9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1359 = 10'h3ca == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1360 = 10'h3cb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1361 = 10'h3cc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1362 = 10'h3cd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1363 = 10'h3ce == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1364 = 10'h3cf == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1365 = 10'h3d0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1366 = 10'h3d1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1367 = 10'h3d2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1368 = 10'h3d3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1369 = 10'h3d4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1370 = 10'h3d5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1371 = 10'h3d6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1372 = 10'h3d7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1373 = 10'h3d8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1374 = 10'h3d9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1375 = 10'h3da == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1376 = 10'h3db == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1377 = 10'h3dc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1378 = 10'h3dd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1379 = 10'h3de == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1380 = 10'h3df == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1381 = 10'h3e0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1382 = 10'h3e1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1383 = 10'h3e2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1384 = 10'h3e3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1385 = 10'h3e4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1386 = 10'h3e5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1387 = 10'h3e6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1388 = 10'h3e7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1389 = 10'h3e8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1390 = 10'h3e9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1391 = 10'h3ea == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1392 = 10'h3eb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1393 = 10'h3ec == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1394 = 10'h3ed == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1395 = 10'h3ee == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1396 = 10'h3ef == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1397 = 10'h3f0 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1398 = 10'h3f1 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1399 = 10'h3f2 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1400 = 10'h3f3 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1401 = 10'h3f4 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1402 = 10'h3f5 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1403 = 10'h3f6 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1404 = 10'h3f7 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1405 = 10'h3f8 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1406 = 10'h3f9 == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1407 = 10'h3fa == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1408 = 10'h3fb == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1409 = 10'h3fc == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1410 = 10'h3fd == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1411 = 10'h3fe == selectedHartReg ? goReg : 1'h0;
  assign _GEN_1412 = 10'h3ff == selectedHartReg ? goReg : 1'h0;
  assign _T_23654 = _T_2863[15:0];
  assign _T_23655 = _T_2863[16];
  assign _T_23656 = _T_2863[17];
  assign _T_23657 = _T_2863[18];
  assign _T_23659 = _T_2863[22:20];
  assign abstractGeneratedI_rd = _T_23685[4:0];
  assign abstractGeneratedS_rs2 = _T_23685[4:0];
  assign _T_23685 = _T_23654 & 16'h1f;
  assign _T_23719 = {abstractGeneratedI_rd,7'h3};
  assign _T_23721 = {17'h7000,_T_23659};
  assign _T_23722 = {_T_23721,_T_23719};
  assign _T_23723 = {_T_23659,5'h0};
  assign _T_23724 = {_T_23723,7'h23};
  assign _T_23725 = {7'h1c,abstractGeneratedS_rs2};
  assign _T_23726 = {_T_23725,5'h0};
  assign _T_23727 = {_T_23726,_T_23724};
  assign _T_23728 = _T_23655 ? _T_23722 : _T_23727;
  assign _T_23733 = _T_23656 ? _T_23728 : 32'h13;
  assign _T_23739 = _T_23657 ? 32'h13 : 32'h100073;
  assign _GEN_2437 = _GEN_5663 ? _T_23733 : abstractGeneratedMem_0;
  assign _GEN_2438 = _GEN_5663 ? _T_23739 : abstractGeneratedMem_1;
  assign _T_23745 = {6'h0,resumeReqRegs_0};
  assign _T_23746 = {_T_23745,_GEN_389};
  assign _T_23748 = {7'h0,_GEN_390};
  assign _T_23750 = {7'h0,_GEN_391};
  assign _T_23752 = {7'h0,_GEN_392};
  assign _T_23754 = {7'h0,_GEN_393};
  assign _T_23756 = {7'h0,_GEN_394};
  assign _T_23758 = {7'h0,_GEN_395};
  assign _T_23760 = {7'h0,_GEN_396};
  assign _T_23762 = {7'h0,_GEN_397};
  assign _T_23764 = {7'h0,_GEN_398};
  assign _T_23766 = {7'h0,_GEN_399};
  assign _T_23768 = {7'h0,_GEN_400};
  assign _T_23770 = {7'h0,_GEN_401};
  assign _T_23772 = {7'h0,_GEN_402};
  assign _T_23774 = {7'h0,_GEN_403};
  assign _T_23776 = {7'h0,_GEN_404};
  assign _T_23778 = {7'h0,_GEN_405};
  assign _T_23780 = {7'h0,_GEN_406};
  assign _T_23782 = {7'h0,_GEN_407};
  assign _T_23784 = {7'h0,_GEN_408};
  assign _T_23786 = {7'h0,_GEN_409};
  assign _T_23788 = {7'h0,_GEN_410};
  assign _T_23790 = {7'h0,_GEN_411};
  assign _T_23792 = {7'h0,_GEN_412};
  assign _T_23794 = {7'h0,_GEN_413};
  assign _T_23796 = {7'h0,_GEN_414};
  assign _T_23798 = {7'h0,_GEN_415};
  assign _T_23800 = {7'h0,_GEN_416};
  assign _T_23802 = {7'h0,_GEN_417};
  assign _T_23804 = {7'h0,_GEN_418};
  assign _T_23806 = {7'h0,_GEN_419};
  assign _T_23808 = {7'h0,_GEN_420};
  assign _T_23810 = {7'h0,_GEN_421};
  assign _T_23812 = {7'h0,_GEN_422};
  assign _T_23814 = {7'h0,_GEN_423};
  assign _T_23816 = {7'h0,_GEN_424};
  assign _T_23818 = {7'h0,_GEN_425};
  assign _T_23820 = {7'h0,_GEN_426};
  assign _T_23822 = {7'h0,_GEN_427};
  assign _T_23824 = {7'h0,_GEN_428};
  assign _T_23826 = {7'h0,_GEN_429};
  assign _T_23828 = {7'h0,_GEN_430};
  assign _T_23830 = {7'h0,_GEN_431};
  assign _T_23832 = {7'h0,_GEN_432};
  assign _T_23834 = {7'h0,_GEN_433};
  assign _T_23836 = {7'h0,_GEN_434};
  assign _T_23838 = {7'h0,_GEN_435};
  assign _T_23840 = {7'h0,_GEN_436};
  assign _T_23842 = {7'h0,_GEN_437};
  assign _T_23844 = {7'h0,_GEN_438};
  assign _T_23846 = {7'h0,_GEN_439};
  assign _T_23848 = {7'h0,_GEN_440};
  assign _T_23850 = {7'h0,_GEN_441};
  assign _T_23852 = {7'h0,_GEN_442};
  assign _T_23854 = {7'h0,_GEN_443};
  assign _T_23856 = {7'h0,_GEN_444};
  assign _T_23858 = {7'h0,_GEN_445};
  assign _T_23860 = {7'h0,_GEN_446};
  assign _T_23862 = {7'h0,_GEN_447};
  assign _T_23864 = {7'h0,_GEN_448};
  assign _T_23866 = {7'h0,_GEN_449};
  assign _T_23868 = {7'h0,_GEN_450};
  assign _T_23870 = {7'h0,_GEN_451};
  assign _T_23872 = {7'h0,_GEN_452};
  assign _T_23874 = {7'h0,_GEN_453};
  assign _T_23876 = {7'h0,_GEN_454};
  assign _T_23878 = {7'h0,_GEN_455};
  assign _T_23880 = {7'h0,_GEN_456};
  assign _T_23882 = {7'h0,_GEN_457};
  assign _T_23884 = {7'h0,_GEN_458};
  assign _T_23886 = {7'h0,_GEN_459};
  assign _T_23888 = {7'h0,_GEN_460};
  assign _T_23890 = {7'h0,_GEN_461};
  assign _T_23892 = {7'h0,_GEN_462};
  assign _T_23894 = {7'h0,_GEN_463};
  assign _T_23896 = {7'h0,_GEN_464};
  assign _T_23898 = {7'h0,_GEN_465};
  assign _T_23900 = {7'h0,_GEN_466};
  assign _T_23902 = {7'h0,_GEN_467};
  assign _T_23904 = {7'h0,_GEN_468};
  assign _T_23906 = {7'h0,_GEN_469};
  assign _T_23908 = {7'h0,_GEN_470};
  assign _T_23910 = {7'h0,_GEN_471};
  assign _T_23912 = {7'h0,_GEN_472};
  assign _T_23914 = {7'h0,_GEN_473};
  assign _T_23916 = {7'h0,_GEN_474};
  assign _T_23918 = {7'h0,_GEN_475};
  assign _T_23920 = {7'h0,_GEN_476};
  assign _T_23922 = {7'h0,_GEN_477};
  assign _T_23924 = {7'h0,_GEN_478};
  assign _T_23926 = {7'h0,_GEN_479};
  assign _T_23928 = {7'h0,_GEN_480};
  assign _T_23930 = {7'h0,_GEN_481};
  assign _T_23932 = {7'h0,_GEN_482};
  assign _T_23934 = {7'h0,_GEN_483};
  assign _T_23936 = {7'h0,_GEN_484};
  assign _T_23938 = {7'h0,_GEN_485};
  assign _T_23940 = {7'h0,_GEN_486};
  assign _T_23942 = {7'h0,_GEN_487};
  assign _T_23944 = {7'h0,_GEN_488};
  assign _T_23946 = {7'h0,_GEN_489};
  assign _T_23948 = {7'h0,_GEN_490};
  assign _T_23950 = {7'h0,_GEN_491};
  assign _T_23952 = {7'h0,_GEN_492};
  assign _T_23954 = {7'h0,_GEN_493};
  assign _T_23956 = {7'h0,_GEN_494};
  assign _T_23958 = {7'h0,_GEN_495};
  assign _T_23960 = {7'h0,_GEN_496};
  assign _T_23962 = {7'h0,_GEN_497};
  assign _T_23964 = {7'h0,_GEN_498};
  assign _T_23966 = {7'h0,_GEN_499};
  assign _T_23968 = {7'h0,_GEN_500};
  assign _T_23970 = {7'h0,_GEN_501};
  assign _T_23972 = {7'h0,_GEN_502};
  assign _T_23974 = {7'h0,_GEN_503};
  assign _T_23976 = {7'h0,_GEN_504};
  assign _T_23978 = {7'h0,_GEN_505};
  assign _T_23980 = {7'h0,_GEN_506};
  assign _T_23982 = {7'h0,_GEN_507};
  assign _T_23984 = {7'h0,_GEN_508};
  assign _T_23986 = {7'h0,_GEN_509};
  assign _T_23988 = {7'h0,_GEN_510};
  assign _T_23990 = {7'h0,_GEN_511};
  assign _T_23992 = {7'h0,_GEN_512};
  assign _T_23994 = {7'h0,_GEN_513};
  assign _T_23996 = {7'h0,_GEN_514};
  assign _T_23998 = {7'h0,_GEN_515};
  assign _T_24000 = {7'h0,_GEN_516};
  assign _T_24002 = {7'h0,_GEN_517};
  assign _T_24004 = {7'h0,_GEN_518};
  assign _T_24006 = {7'h0,_GEN_519};
  assign _T_24008 = {7'h0,_GEN_520};
  assign _T_24010 = {7'h0,_GEN_521};
  assign _T_24012 = {7'h0,_GEN_522};
  assign _T_24014 = {7'h0,_GEN_523};
  assign _T_24016 = {7'h0,_GEN_524};
  assign _T_24018 = {7'h0,_GEN_525};
  assign _T_24020 = {7'h0,_GEN_526};
  assign _T_24022 = {7'h0,_GEN_527};
  assign _T_24024 = {7'h0,_GEN_528};
  assign _T_24026 = {7'h0,_GEN_529};
  assign _T_24028 = {7'h0,_GEN_530};
  assign _T_24030 = {7'h0,_GEN_531};
  assign _T_24032 = {7'h0,_GEN_532};
  assign _T_24034 = {7'h0,_GEN_533};
  assign _T_24036 = {7'h0,_GEN_534};
  assign _T_24038 = {7'h0,_GEN_535};
  assign _T_24040 = {7'h0,_GEN_536};
  assign _T_24042 = {7'h0,_GEN_537};
  assign _T_24044 = {7'h0,_GEN_538};
  assign _T_24046 = {7'h0,_GEN_539};
  assign _T_24048 = {7'h0,_GEN_540};
  assign _T_24050 = {7'h0,_GEN_541};
  assign _T_24052 = {7'h0,_GEN_542};
  assign _T_24054 = {7'h0,_GEN_543};
  assign _T_24056 = {7'h0,_GEN_544};
  assign _T_24058 = {7'h0,_GEN_545};
  assign _T_24060 = {7'h0,_GEN_546};
  assign _T_24062 = {7'h0,_GEN_547};
  assign _T_24064 = {7'h0,_GEN_548};
  assign _T_24066 = {7'h0,_GEN_549};
  assign _T_24068 = {7'h0,_GEN_550};
  assign _T_24070 = {7'h0,_GEN_551};
  assign _T_24072 = {7'h0,_GEN_552};
  assign _T_24074 = {7'h0,_GEN_553};
  assign _T_24076 = {7'h0,_GEN_554};
  assign _T_24078 = {7'h0,_GEN_555};
  assign _T_24080 = {7'h0,_GEN_556};
  assign _T_24082 = {7'h0,_GEN_557};
  assign _T_24084 = {7'h0,_GEN_558};
  assign _T_24086 = {7'h0,_GEN_559};
  assign _T_24088 = {7'h0,_GEN_560};
  assign _T_24090 = {7'h0,_GEN_561};
  assign _T_24092 = {7'h0,_GEN_562};
  assign _T_24094 = {7'h0,_GEN_563};
  assign _T_24096 = {7'h0,_GEN_564};
  assign _T_24098 = {7'h0,_GEN_565};
  assign _T_24100 = {7'h0,_GEN_566};
  assign _T_24102 = {7'h0,_GEN_567};
  assign _T_24104 = {7'h0,_GEN_568};
  assign _T_24106 = {7'h0,_GEN_569};
  assign _T_24108 = {7'h0,_GEN_570};
  assign _T_24110 = {7'h0,_GEN_571};
  assign _T_24112 = {7'h0,_GEN_572};
  assign _T_24114 = {7'h0,_GEN_573};
  assign _T_24116 = {7'h0,_GEN_574};
  assign _T_24118 = {7'h0,_GEN_575};
  assign _T_24120 = {7'h0,_GEN_576};
  assign _T_24122 = {7'h0,_GEN_577};
  assign _T_24124 = {7'h0,_GEN_578};
  assign _T_24126 = {7'h0,_GEN_579};
  assign _T_24128 = {7'h0,_GEN_580};
  assign _T_24130 = {7'h0,_GEN_581};
  assign _T_24132 = {7'h0,_GEN_582};
  assign _T_24134 = {7'h0,_GEN_583};
  assign _T_24136 = {7'h0,_GEN_584};
  assign _T_24138 = {7'h0,_GEN_585};
  assign _T_24140 = {7'h0,_GEN_586};
  assign _T_24142 = {7'h0,_GEN_587};
  assign _T_24144 = {7'h0,_GEN_588};
  assign _T_24146 = {7'h0,_GEN_589};
  assign _T_24148 = {7'h0,_GEN_590};
  assign _T_24150 = {7'h0,_GEN_591};
  assign _T_24152 = {7'h0,_GEN_592};
  assign _T_24154 = {7'h0,_GEN_593};
  assign _T_24156 = {7'h0,_GEN_594};
  assign _T_24158 = {7'h0,_GEN_595};
  assign _T_24160 = {7'h0,_GEN_596};
  assign _T_24162 = {7'h0,_GEN_597};
  assign _T_24164 = {7'h0,_GEN_598};
  assign _T_24166 = {7'h0,_GEN_599};
  assign _T_24168 = {7'h0,_GEN_600};
  assign _T_24170 = {7'h0,_GEN_601};
  assign _T_24172 = {7'h0,_GEN_602};
  assign _T_24174 = {7'h0,_GEN_603};
  assign _T_24176 = {7'h0,_GEN_604};
  assign _T_24178 = {7'h0,_GEN_605};
  assign _T_24180 = {7'h0,_GEN_606};
  assign _T_24182 = {7'h0,_GEN_607};
  assign _T_24184 = {7'h0,_GEN_608};
  assign _T_24186 = {7'h0,_GEN_609};
  assign _T_24188 = {7'h0,_GEN_610};
  assign _T_24190 = {7'h0,_GEN_611};
  assign _T_24192 = {7'h0,_GEN_612};
  assign _T_24194 = {7'h0,_GEN_613};
  assign _T_24196 = {7'h0,_GEN_614};
  assign _T_24198 = {7'h0,_GEN_615};
  assign _T_24200 = {7'h0,_GEN_616};
  assign _T_24202 = {7'h0,_GEN_617};
  assign _T_24204 = {7'h0,_GEN_618};
  assign _T_24206 = {7'h0,_GEN_619};
  assign _T_24208 = {7'h0,_GEN_620};
  assign _T_24210 = {7'h0,_GEN_621};
  assign _T_24212 = {7'h0,_GEN_622};
  assign _T_24214 = {7'h0,_GEN_623};
  assign _T_24216 = {7'h0,_GEN_624};
  assign _T_24218 = {7'h0,_GEN_625};
  assign _T_24220 = {7'h0,_GEN_626};
  assign _T_24222 = {7'h0,_GEN_627};
  assign _T_24224 = {7'h0,_GEN_628};
  assign _T_24226 = {7'h0,_GEN_629};
  assign _T_24228 = {7'h0,_GEN_630};
  assign _T_24230 = {7'h0,_GEN_631};
  assign _T_24232 = {7'h0,_GEN_632};
  assign _T_24234 = {7'h0,_GEN_633};
  assign _T_24236 = {7'h0,_GEN_634};
  assign _T_24238 = {7'h0,_GEN_635};
  assign _T_24240 = {7'h0,_GEN_636};
  assign _T_24242 = {7'h0,_GEN_637};
  assign _T_24244 = {7'h0,_GEN_638};
  assign _T_24246 = {7'h0,_GEN_639};
  assign _T_24248 = {7'h0,_GEN_640};
  assign _T_24250 = {7'h0,_GEN_641};
  assign _T_24252 = {7'h0,_GEN_642};
  assign _T_24254 = {7'h0,_GEN_643};
  assign _T_24256 = {7'h0,_GEN_644};
  assign _T_24258 = {7'h0,_GEN_645};
  assign _T_24260 = {7'h0,_GEN_646};
  assign _T_24262 = {7'h0,_GEN_647};
  assign _T_24264 = {7'h0,_GEN_648};
  assign _T_24266 = {7'h0,_GEN_649};
  assign _T_24268 = {7'h0,_GEN_650};
  assign _T_24270 = {7'h0,_GEN_651};
  assign _T_24272 = {7'h0,_GEN_652};
  assign _T_24274 = {7'h0,_GEN_653};
  assign _T_24276 = {7'h0,_GEN_654};
  assign _T_24278 = {7'h0,_GEN_655};
  assign _T_24280 = {7'h0,_GEN_656};
  assign _T_24282 = {7'h0,_GEN_657};
  assign _T_24284 = {7'h0,_GEN_658};
  assign _T_24286 = {7'h0,_GEN_659};
  assign _T_24288 = {7'h0,_GEN_660};
  assign _T_24290 = {7'h0,_GEN_661};
  assign _T_24292 = {7'h0,_GEN_662};
  assign _T_24294 = {7'h0,_GEN_663};
  assign _T_24296 = {7'h0,_GEN_664};
  assign _T_24298 = {7'h0,_GEN_665};
  assign _T_24300 = {7'h0,_GEN_666};
  assign _T_24302 = {7'h0,_GEN_667};
  assign _T_24304 = {7'h0,_GEN_668};
  assign _T_24306 = {7'h0,_GEN_669};
  assign _T_24308 = {7'h0,_GEN_670};
  assign _T_24310 = {7'h0,_GEN_671};
  assign _T_24312 = {7'h0,_GEN_672};
  assign _T_24314 = {7'h0,_GEN_673};
  assign _T_24316 = {7'h0,_GEN_674};
  assign _T_24318 = {7'h0,_GEN_675};
  assign _T_24320 = {7'h0,_GEN_676};
  assign _T_24322 = {7'h0,_GEN_677};
  assign _T_24324 = {7'h0,_GEN_678};
  assign _T_24326 = {7'h0,_GEN_679};
  assign _T_24328 = {7'h0,_GEN_680};
  assign _T_24330 = {7'h0,_GEN_681};
  assign _T_24332 = {7'h0,_GEN_682};
  assign _T_24334 = {7'h0,_GEN_683};
  assign _T_24336 = {7'h0,_GEN_684};
  assign _T_24338 = {7'h0,_GEN_685};
  assign _T_24340 = {7'h0,_GEN_686};
  assign _T_24342 = {7'h0,_GEN_687};
  assign _T_24344 = {7'h0,_GEN_688};
  assign _T_24346 = {7'h0,_GEN_689};
  assign _T_24348 = {7'h0,_GEN_690};
  assign _T_24350 = {7'h0,_GEN_691};
  assign _T_24352 = {7'h0,_GEN_692};
  assign _T_24354 = {7'h0,_GEN_693};
  assign _T_24356 = {7'h0,_GEN_694};
  assign _T_24358 = {7'h0,_GEN_695};
  assign _T_24360 = {7'h0,_GEN_696};
  assign _T_24362 = {7'h0,_GEN_697};
  assign _T_24364 = {7'h0,_GEN_698};
  assign _T_24366 = {7'h0,_GEN_699};
  assign _T_24368 = {7'h0,_GEN_700};
  assign _T_24370 = {7'h0,_GEN_701};
  assign _T_24372 = {7'h0,_GEN_702};
  assign _T_24374 = {7'h0,_GEN_703};
  assign _T_24376 = {7'h0,_GEN_704};
  assign _T_24378 = {7'h0,_GEN_705};
  assign _T_24380 = {7'h0,_GEN_706};
  assign _T_24382 = {7'h0,_GEN_707};
  assign _T_24384 = {7'h0,_GEN_708};
  assign _T_24386 = {7'h0,_GEN_709};
  assign _T_24388 = {7'h0,_GEN_710};
  assign _T_24390 = {7'h0,_GEN_711};
  assign _T_24392 = {7'h0,_GEN_712};
  assign _T_24394 = {7'h0,_GEN_713};
  assign _T_24396 = {7'h0,_GEN_714};
  assign _T_24398 = {7'h0,_GEN_715};
  assign _T_24400 = {7'h0,_GEN_716};
  assign _T_24402 = {7'h0,_GEN_717};
  assign _T_24404 = {7'h0,_GEN_718};
  assign _T_24406 = {7'h0,_GEN_719};
  assign _T_24408 = {7'h0,_GEN_720};
  assign _T_24410 = {7'h0,_GEN_721};
  assign _T_24412 = {7'h0,_GEN_722};
  assign _T_24414 = {7'h0,_GEN_723};
  assign _T_24416 = {7'h0,_GEN_724};
  assign _T_24418 = {7'h0,_GEN_725};
  assign _T_24420 = {7'h0,_GEN_726};
  assign _T_24422 = {7'h0,_GEN_727};
  assign _T_24424 = {7'h0,_GEN_728};
  assign _T_24426 = {7'h0,_GEN_729};
  assign _T_24428 = {7'h0,_GEN_730};
  assign _T_24430 = {7'h0,_GEN_731};
  assign _T_24432 = {7'h0,_GEN_732};
  assign _T_24434 = {7'h0,_GEN_733};
  assign _T_24436 = {7'h0,_GEN_734};
  assign _T_24438 = {7'h0,_GEN_735};
  assign _T_24440 = {7'h0,_GEN_736};
  assign _T_24442 = {7'h0,_GEN_737};
  assign _T_24444 = {7'h0,_GEN_738};
  assign _T_24446 = {7'h0,_GEN_739};
  assign _T_24448 = {7'h0,_GEN_740};
  assign _T_24450 = {7'h0,_GEN_741};
  assign _T_24452 = {7'h0,_GEN_742};
  assign _T_24454 = {7'h0,_GEN_743};
  assign _T_24456 = {7'h0,_GEN_744};
  assign _T_24458 = {7'h0,_GEN_745};
  assign _T_24460 = {7'h0,_GEN_746};
  assign _T_24462 = {7'h0,_GEN_747};
  assign _T_24464 = {7'h0,_GEN_748};
  assign _T_24466 = {7'h0,_GEN_749};
  assign _T_24468 = {7'h0,_GEN_750};
  assign _T_24470 = {7'h0,_GEN_751};
  assign _T_24472 = {7'h0,_GEN_752};
  assign _T_24474 = {7'h0,_GEN_753};
  assign _T_24476 = {7'h0,_GEN_754};
  assign _T_24478 = {7'h0,_GEN_755};
  assign _T_24480 = {7'h0,_GEN_756};
  assign _T_24482 = {7'h0,_GEN_757};
  assign _T_24484 = {7'h0,_GEN_758};
  assign _T_24486 = {7'h0,_GEN_759};
  assign _T_24488 = {7'h0,_GEN_760};
  assign _T_24490 = {7'h0,_GEN_761};
  assign _T_24492 = {7'h0,_GEN_762};
  assign _T_24494 = {7'h0,_GEN_763};
  assign _T_24496 = {7'h0,_GEN_764};
  assign _T_24498 = {7'h0,_GEN_765};
  assign _T_24500 = {7'h0,_GEN_766};
  assign _T_24502 = {7'h0,_GEN_767};
  assign _T_24504 = {7'h0,_GEN_768};
  assign _T_24506 = {7'h0,_GEN_769};
  assign _T_24508 = {7'h0,_GEN_770};
  assign _T_24510 = {7'h0,_GEN_771};
  assign _T_24512 = {7'h0,_GEN_772};
  assign _T_24514 = {7'h0,_GEN_773};
  assign _T_24516 = {7'h0,_GEN_774};
  assign _T_24518 = {7'h0,_GEN_775};
  assign _T_24520 = {7'h0,_GEN_776};
  assign _T_24522 = {7'h0,_GEN_777};
  assign _T_24524 = {7'h0,_GEN_778};
  assign _T_24526 = {7'h0,_GEN_779};
  assign _T_24528 = {7'h0,_GEN_780};
  assign _T_24530 = {7'h0,_GEN_781};
  assign _T_24532 = {7'h0,_GEN_782};
  assign _T_24534 = {7'h0,_GEN_783};
  assign _T_24536 = {7'h0,_GEN_784};
  assign _T_24538 = {7'h0,_GEN_785};
  assign _T_24540 = {7'h0,_GEN_786};
  assign _T_24542 = {7'h0,_GEN_787};
  assign _T_24544 = {7'h0,_GEN_788};
  assign _T_24546 = {7'h0,_GEN_789};
  assign _T_24548 = {7'h0,_GEN_790};
  assign _T_24550 = {7'h0,_GEN_791};
  assign _T_24552 = {7'h0,_GEN_792};
  assign _T_24554 = {7'h0,_GEN_793};
  assign _T_24556 = {7'h0,_GEN_794};
  assign _T_24558 = {7'h0,_GEN_795};
  assign _T_24560 = {7'h0,_GEN_796};
  assign _T_24562 = {7'h0,_GEN_797};
  assign _T_24564 = {7'h0,_GEN_798};
  assign _T_24566 = {7'h0,_GEN_799};
  assign _T_24568 = {7'h0,_GEN_800};
  assign _T_24570 = {7'h0,_GEN_801};
  assign _T_24572 = {7'h0,_GEN_802};
  assign _T_24574 = {7'h0,_GEN_803};
  assign _T_24576 = {7'h0,_GEN_804};
  assign _T_24578 = {7'h0,_GEN_805};
  assign _T_24580 = {7'h0,_GEN_806};
  assign _T_24582 = {7'h0,_GEN_807};
  assign _T_24584 = {7'h0,_GEN_808};
  assign _T_24586 = {7'h0,_GEN_809};
  assign _T_24588 = {7'h0,_GEN_810};
  assign _T_24590 = {7'h0,_GEN_811};
  assign _T_24592 = {7'h0,_GEN_812};
  assign _T_24594 = {7'h0,_GEN_813};
  assign _T_24596 = {7'h0,_GEN_814};
  assign _T_24598 = {7'h0,_GEN_815};
  assign _T_24600 = {7'h0,_GEN_816};
  assign _T_24602 = {7'h0,_GEN_817};
  assign _T_24604 = {7'h0,_GEN_818};
  assign _T_24606 = {7'h0,_GEN_819};
  assign _T_24608 = {7'h0,_GEN_820};
  assign _T_24610 = {7'h0,_GEN_821};
  assign _T_24612 = {7'h0,_GEN_822};
  assign _T_24614 = {7'h0,_GEN_823};
  assign _T_24616 = {7'h0,_GEN_824};
  assign _T_24618 = {7'h0,_GEN_825};
  assign _T_24620 = {7'h0,_GEN_826};
  assign _T_24622 = {7'h0,_GEN_827};
  assign _T_24624 = {7'h0,_GEN_828};
  assign _T_24626 = {7'h0,_GEN_829};
  assign _T_24628 = {7'h0,_GEN_830};
  assign _T_24630 = {7'h0,_GEN_831};
  assign _T_24632 = {7'h0,_GEN_832};
  assign _T_24634 = {7'h0,_GEN_833};
  assign _T_24636 = {7'h0,_GEN_834};
  assign _T_24638 = {7'h0,_GEN_835};
  assign _T_24640 = {7'h0,_GEN_836};
  assign _T_24642 = {7'h0,_GEN_837};
  assign _T_24644 = {7'h0,_GEN_838};
  assign _T_24646 = {7'h0,_GEN_839};
  assign _T_24648 = {7'h0,_GEN_840};
  assign _T_24650 = {7'h0,_GEN_841};
  assign _T_24652 = {7'h0,_GEN_842};
  assign _T_24654 = {7'h0,_GEN_843};
  assign _T_24656 = {7'h0,_GEN_844};
  assign _T_24658 = {7'h0,_GEN_845};
  assign _T_24660 = {7'h0,_GEN_846};
  assign _T_24662 = {7'h0,_GEN_847};
  assign _T_24664 = {7'h0,_GEN_848};
  assign _T_24666 = {7'h0,_GEN_849};
  assign _T_24668 = {7'h0,_GEN_850};
  assign _T_24670 = {7'h0,_GEN_851};
  assign _T_24672 = {7'h0,_GEN_852};
  assign _T_24674 = {7'h0,_GEN_853};
  assign _T_24676 = {7'h0,_GEN_854};
  assign _T_24678 = {7'h0,_GEN_855};
  assign _T_24680 = {7'h0,_GEN_856};
  assign _T_24682 = {7'h0,_GEN_857};
  assign _T_24684 = {7'h0,_GEN_858};
  assign _T_24686 = {7'h0,_GEN_859};
  assign _T_24688 = {7'h0,_GEN_860};
  assign _T_24690 = {7'h0,_GEN_861};
  assign _T_24692 = {7'h0,_GEN_862};
  assign _T_24694 = {7'h0,_GEN_863};
  assign _T_24696 = {7'h0,_GEN_864};
  assign _T_24698 = {7'h0,_GEN_865};
  assign _T_24700 = {7'h0,_GEN_866};
  assign _T_24702 = {7'h0,_GEN_867};
  assign _T_24704 = {7'h0,_GEN_868};
  assign _T_24706 = {7'h0,_GEN_869};
  assign _T_24708 = {7'h0,_GEN_870};
  assign _T_24710 = {7'h0,_GEN_871};
  assign _T_24712 = {7'h0,_GEN_872};
  assign _T_24714 = {7'h0,_GEN_873};
  assign _T_24716 = {7'h0,_GEN_874};
  assign _T_24718 = {7'h0,_GEN_875};
  assign _T_24720 = {7'h0,_GEN_876};
  assign _T_24722 = {7'h0,_GEN_877};
  assign _T_24724 = {7'h0,_GEN_878};
  assign _T_24726 = {7'h0,_GEN_879};
  assign _T_24728 = {7'h0,_GEN_880};
  assign _T_24730 = {7'h0,_GEN_881};
  assign _T_24732 = {7'h0,_GEN_882};
  assign _T_24734 = {7'h0,_GEN_883};
  assign _T_24736 = {7'h0,_GEN_884};
  assign _T_24738 = {7'h0,_GEN_885};
  assign _T_24740 = {7'h0,_GEN_886};
  assign _T_24742 = {7'h0,_GEN_887};
  assign _T_24744 = {7'h0,_GEN_888};
  assign _T_24746 = {7'h0,_GEN_889};
  assign _T_24748 = {7'h0,_GEN_890};
  assign _T_24750 = {7'h0,_GEN_891};
  assign _T_24752 = {7'h0,_GEN_892};
  assign _T_24754 = {7'h0,_GEN_893};
  assign _T_24756 = {7'h0,_GEN_894};
  assign _T_24758 = {7'h0,_GEN_895};
  assign _T_24760 = {7'h0,_GEN_896};
  assign _T_24762 = {7'h0,_GEN_897};
  assign _T_24764 = {7'h0,_GEN_898};
  assign _T_24766 = {7'h0,_GEN_899};
  assign _T_24768 = {7'h0,_GEN_900};
  assign _T_24770 = {7'h0,_GEN_901};
  assign _T_24772 = {7'h0,_GEN_902};
  assign _T_24774 = {7'h0,_GEN_903};
  assign _T_24776 = {7'h0,_GEN_904};
  assign _T_24778 = {7'h0,_GEN_905};
  assign _T_24780 = {7'h0,_GEN_906};
  assign _T_24782 = {7'h0,_GEN_907};
  assign _T_24784 = {7'h0,_GEN_908};
  assign _T_24786 = {7'h0,_GEN_909};
  assign _T_24788 = {7'h0,_GEN_910};
  assign _T_24790 = {7'h0,_GEN_911};
  assign _T_24792 = {7'h0,_GEN_912};
  assign _T_24794 = {7'h0,_GEN_913};
  assign _T_24796 = {7'h0,_GEN_914};
  assign _T_24798 = {7'h0,_GEN_915};
  assign _T_24800 = {7'h0,_GEN_916};
  assign _T_24802 = {7'h0,_GEN_917};
  assign _T_24804 = {7'h0,_GEN_918};
  assign _T_24806 = {7'h0,_GEN_919};
  assign _T_24808 = {7'h0,_GEN_920};
  assign _T_24810 = {7'h0,_GEN_921};
  assign _T_24812 = {7'h0,_GEN_922};
  assign _T_24814 = {7'h0,_GEN_923};
  assign _T_24816 = {7'h0,_GEN_924};
  assign _T_24818 = {7'h0,_GEN_925};
  assign _T_24820 = {7'h0,_GEN_926};
  assign _T_24822 = {7'h0,_GEN_927};
  assign _T_24824 = {7'h0,_GEN_928};
  assign _T_24826 = {7'h0,_GEN_929};
  assign _T_24828 = {7'h0,_GEN_930};
  assign _T_24830 = {7'h0,_GEN_931};
  assign _T_24832 = {7'h0,_GEN_932};
  assign _T_24834 = {7'h0,_GEN_933};
  assign _T_24836 = {7'h0,_GEN_934};
  assign _T_24838 = {7'h0,_GEN_935};
  assign _T_24840 = {7'h0,_GEN_936};
  assign _T_24842 = {7'h0,_GEN_937};
  assign _T_24844 = {7'h0,_GEN_938};
  assign _T_24846 = {7'h0,_GEN_939};
  assign _T_24848 = {7'h0,_GEN_940};
  assign _T_24850 = {7'h0,_GEN_941};
  assign _T_24852 = {7'h0,_GEN_942};
  assign _T_24854 = {7'h0,_GEN_943};
  assign _T_24856 = {7'h0,_GEN_944};
  assign _T_24858 = {7'h0,_GEN_945};
  assign _T_24860 = {7'h0,_GEN_946};
  assign _T_24862 = {7'h0,_GEN_947};
  assign _T_24864 = {7'h0,_GEN_948};
  assign _T_24866 = {7'h0,_GEN_949};
  assign _T_24868 = {7'h0,_GEN_950};
  assign _T_24870 = {7'h0,_GEN_951};
  assign _T_24872 = {7'h0,_GEN_952};
  assign _T_24874 = {7'h0,_GEN_953};
  assign _T_24876 = {7'h0,_GEN_954};
  assign _T_24878 = {7'h0,_GEN_955};
  assign _T_24880 = {7'h0,_GEN_956};
  assign _T_24882 = {7'h0,_GEN_957};
  assign _T_24884 = {7'h0,_GEN_958};
  assign _T_24886 = {7'h0,_GEN_959};
  assign _T_24888 = {7'h0,_GEN_960};
  assign _T_24890 = {7'h0,_GEN_961};
  assign _T_24892 = {7'h0,_GEN_962};
  assign _T_24894 = {7'h0,_GEN_963};
  assign _T_24896 = {7'h0,_GEN_964};
  assign _T_24898 = {7'h0,_GEN_965};
  assign _T_24900 = {7'h0,_GEN_966};
  assign _T_24902 = {7'h0,_GEN_967};
  assign _T_24904 = {7'h0,_GEN_968};
  assign _T_24906 = {7'h0,_GEN_969};
  assign _T_24908 = {7'h0,_GEN_970};
  assign _T_24910 = {7'h0,_GEN_971};
  assign _T_24912 = {7'h0,_GEN_972};
  assign _T_24914 = {7'h0,_GEN_973};
  assign _T_24916 = {7'h0,_GEN_974};
  assign _T_24918 = {7'h0,_GEN_975};
  assign _T_24920 = {7'h0,_GEN_976};
  assign _T_24922 = {7'h0,_GEN_977};
  assign _T_24924 = {7'h0,_GEN_978};
  assign _T_24926 = {7'h0,_GEN_979};
  assign _T_24928 = {7'h0,_GEN_980};
  assign _T_24930 = {7'h0,_GEN_981};
  assign _T_24932 = {7'h0,_GEN_982};
  assign _T_24934 = {7'h0,_GEN_983};
  assign _T_24936 = {7'h0,_GEN_984};
  assign _T_24938 = {7'h0,_GEN_985};
  assign _T_24940 = {7'h0,_GEN_986};
  assign _T_24942 = {7'h0,_GEN_987};
  assign _T_24944 = {7'h0,_GEN_988};
  assign _T_24946 = {7'h0,_GEN_989};
  assign _T_24948 = {7'h0,_GEN_990};
  assign _T_24950 = {7'h0,_GEN_991};
  assign _T_24952 = {7'h0,_GEN_992};
  assign _T_24954 = {7'h0,_GEN_993};
  assign _T_24956 = {7'h0,_GEN_994};
  assign _T_24958 = {7'h0,_GEN_995};
  assign _T_24960 = {7'h0,_GEN_996};
  assign _T_24962 = {7'h0,_GEN_997};
  assign _T_24964 = {7'h0,_GEN_998};
  assign _T_24966 = {7'h0,_GEN_999};
  assign _T_24968 = {7'h0,_GEN_1000};
  assign _T_24970 = {7'h0,_GEN_1001};
  assign _T_24972 = {7'h0,_GEN_1002};
  assign _T_24974 = {7'h0,_GEN_1003};
  assign _T_24976 = {7'h0,_GEN_1004};
  assign _T_24978 = {7'h0,_GEN_1005};
  assign _T_24980 = {7'h0,_GEN_1006};
  assign _T_24982 = {7'h0,_GEN_1007};
  assign _T_24984 = {7'h0,_GEN_1008};
  assign _T_24986 = {7'h0,_GEN_1009};
  assign _T_24988 = {7'h0,_GEN_1010};
  assign _T_24990 = {7'h0,_GEN_1011};
  assign _T_24992 = {7'h0,_GEN_1012};
  assign _T_24994 = {7'h0,_GEN_1013};
  assign _T_24996 = {7'h0,_GEN_1014};
  assign _T_24998 = {7'h0,_GEN_1015};
  assign _T_25000 = {7'h0,_GEN_1016};
  assign _T_25002 = {7'h0,_GEN_1017};
  assign _T_25004 = {7'h0,_GEN_1018};
  assign _T_25006 = {7'h0,_GEN_1019};
  assign _T_25008 = {7'h0,_GEN_1020};
  assign _T_25010 = {7'h0,_GEN_1021};
  assign _T_25012 = {7'h0,_GEN_1022};
  assign _T_25014 = {7'h0,_GEN_1023};
  assign _T_25016 = {7'h0,_GEN_1024};
  assign _T_25018 = {7'h0,_GEN_1025};
  assign _T_25020 = {7'h0,_GEN_1026};
  assign _T_25022 = {7'h0,_GEN_1027};
  assign _T_25024 = {7'h0,_GEN_1028};
  assign _T_25026 = {7'h0,_GEN_1029};
  assign _T_25028 = {7'h0,_GEN_1030};
  assign _T_25030 = {7'h0,_GEN_1031};
  assign _T_25032 = {7'h0,_GEN_1032};
  assign _T_25034 = {7'h0,_GEN_1033};
  assign _T_25036 = {7'h0,_GEN_1034};
  assign _T_25038 = {7'h0,_GEN_1035};
  assign _T_25040 = {7'h0,_GEN_1036};
  assign _T_25042 = {7'h0,_GEN_1037};
  assign _T_25044 = {7'h0,_GEN_1038};
  assign _T_25046 = {7'h0,_GEN_1039};
  assign _T_25048 = {7'h0,_GEN_1040};
  assign _T_25050 = {7'h0,_GEN_1041};
  assign _T_25052 = {7'h0,_GEN_1042};
  assign _T_25054 = {7'h0,_GEN_1043};
  assign _T_25056 = {7'h0,_GEN_1044};
  assign _T_25058 = {7'h0,_GEN_1045};
  assign _T_25060 = {7'h0,_GEN_1046};
  assign _T_25062 = {7'h0,_GEN_1047};
  assign _T_25064 = {7'h0,_GEN_1048};
  assign _T_25066 = {7'h0,_GEN_1049};
  assign _T_25068 = {7'h0,_GEN_1050};
  assign _T_25070 = {7'h0,_GEN_1051};
  assign _T_25072 = {7'h0,_GEN_1052};
  assign _T_25074 = {7'h0,_GEN_1053};
  assign _T_25076 = {7'h0,_GEN_1054};
  assign _T_25078 = {7'h0,_GEN_1055};
  assign _T_25080 = {7'h0,_GEN_1056};
  assign _T_25082 = {7'h0,_GEN_1057};
  assign _T_25084 = {7'h0,_GEN_1058};
  assign _T_25086 = {7'h0,_GEN_1059};
  assign _T_25088 = {7'h0,_GEN_1060};
  assign _T_25090 = {7'h0,_GEN_1061};
  assign _T_25092 = {7'h0,_GEN_1062};
  assign _T_25094 = {7'h0,_GEN_1063};
  assign _T_25096 = {7'h0,_GEN_1064};
  assign _T_25098 = {7'h0,_GEN_1065};
  assign _T_25100 = {7'h0,_GEN_1066};
  assign _T_25102 = {7'h0,_GEN_1067};
  assign _T_25104 = {7'h0,_GEN_1068};
  assign _T_25106 = {7'h0,_GEN_1069};
  assign _T_25108 = {7'h0,_GEN_1070};
  assign _T_25110 = {7'h0,_GEN_1071};
  assign _T_25112 = {7'h0,_GEN_1072};
  assign _T_25114 = {7'h0,_GEN_1073};
  assign _T_25116 = {7'h0,_GEN_1074};
  assign _T_25118 = {7'h0,_GEN_1075};
  assign _T_25120 = {7'h0,_GEN_1076};
  assign _T_25122 = {7'h0,_GEN_1077};
  assign _T_25124 = {7'h0,_GEN_1078};
  assign _T_25126 = {7'h0,_GEN_1079};
  assign _T_25128 = {7'h0,_GEN_1080};
  assign _T_25130 = {7'h0,_GEN_1081};
  assign _T_25132 = {7'h0,_GEN_1082};
  assign _T_25134 = {7'h0,_GEN_1083};
  assign _T_25136 = {7'h0,_GEN_1084};
  assign _T_25138 = {7'h0,_GEN_1085};
  assign _T_25140 = {7'h0,_GEN_1086};
  assign _T_25142 = {7'h0,_GEN_1087};
  assign _T_25144 = {7'h0,_GEN_1088};
  assign _T_25146 = {7'h0,_GEN_1089};
  assign _T_25148 = {7'h0,_GEN_1090};
  assign _T_25150 = {7'h0,_GEN_1091};
  assign _T_25152 = {7'h0,_GEN_1092};
  assign _T_25154 = {7'h0,_GEN_1093};
  assign _T_25156 = {7'h0,_GEN_1094};
  assign _T_25158 = {7'h0,_GEN_1095};
  assign _T_25160 = {7'h0,_GEN_1096};
  assign _T_25162 = {7'h0,_GEN_1097};
  assign _T_25164 = {7'h0,_GEN_1098};
  assign _T_25166 = {7'h0,_GEN_1099};
  assign _T_25168 = {7'h0,_GEN_1100};
  assign _T_25170 = {7'h0,_GEN_1101};
  assign _T_25172 = {7'h0,_GEN_1102};
  assign _T_25174 = {7'h0,_GEN_1103};
  assign _T_25176 = {7'h0,_GEN_1104};
  assign _T_25178 = {7'h0,_GEN_1105};
  assign _T_25180 = {7'h0,_GEN_1106};
  assign _T_25182 = {7'h0,_GEN_1107};
  assign _T_25184 = {7'h0,_GEN_1108};
  assign _T_25186 = {7'h0,_GEN_1109};
  assign _T_25188 = {7'h0,_GEN_1110};
  assign _T_25190 = {7'h0,_GEN_1111};
  assign _T_25192 = {7'h0,_GEN_1112};
  assign _T_25194 = {7'h0,_GEN_1113};
  assign _T_25196 = {7'h0,_GEN_1114};
  assign _T_25198 = {7'h0,_GEN_1115};
  assign _T_25200 = {7'h0,_GEN_1116};
  assign _T_25202 = {7'h0,_GEN_1117};
  assign _T_25204 = {7'h0,_GEN_1118};
  assign _T_25206 = {7'h0,_GEN_1119};
  assign _T_25208 = {7'h0,_GEN_1120};
  assign _T_25210 = {7'h0,_GEN_1121};
  assign _T_25212 = {7'h0,_GEN_1122};
  assign _T_25214 = {7'h0,_GEN_1123};
  assign _T_25216 = {7'h0,_GEN_1124};
  assign _T_25218 = {7'h0,_GEN_1125};
  assign _T_25220 = {7'h0,_GEN_1126};
  assign _T_25222 = {7'h0,_GEN_1127};
  assign _T_25224 = {7'h0,_GEN_1128};
  assign _T_25226 = {7'h0,_GEN_1129};
  assign _T_25228 = {7'h0,_GEN_1130};
  assign _T_25230 = {7'h0,_GEN_1131};
  assign _T_25232 = {7'h0,_GEN_1132};
  assign _T_25234 = {7'h0,_GEN_1133};
  assign _T_25236 = {7'h0,_GEN_1134};
  assign _T_25238 = {7'h0,_GEN_1135};
  assign _T_25240 = {7'h0,_GEN_1136};
  assign _T_25242 = {7'h0,_GEN_1137};
  assign _T_25244 = {7'h0,_GEN_1138};
  assign _T_25246 = {7'h0,_GEN_1139};
  assign _T_25248 = {7'h0,_GEN_1140};
  assign _T_25250 = {7'h0,_GEN_1141};
  assign _T_25252 = {7'h0,_GEN_1142};
  assign _T_25254 = {7'h0,_GEN_1143};
  assign _T_25256 = {7'h0,_GEN_1144};
  assign _T_25258 = {7'h0,_GEN_1145};
  assign _T_25260 = {7'h0,_GEN_1146};
  assign _T_25262 = {7'h0,_GEN_1147};
  assign _T_25264 = {7'h0,_GEN_1148};
  assign _T_25266 = {7'h0,_GEN_1149};
  assign _T_25268 = {7'h0,_GEN_1150};
  assign _T_25270 = {7'h0,_GEN_1151};
  assign _T_25272 = {7'h0,_GEN_1152};
  assign _T_25274 = {7'h0,_GEN_1153};
  assign _T_25276 = {7'h0,_GEN_1154};
  assign _T_25278 = {7'h0,_GEN_1155};
  assign _T_25280 = {7'h0,_GEN_1156};
  assign _T_25282 = {7'h0,_GEN_1157};
  assign _T_25284 = {7'h0,_GEN_1158};
  assign _T_25286 = {7'h0,_GEN_1159};
  assign _T_25288 = {7'h0,_GEN_1160};
  assign _T_25290 = {7'h0,_GEN_1161};
  assign _T_25292 = {7'h0,_GEN_1162};
  assign _T_25294 = {7'h0,_GEN_1163};
  assign _T_25296 = {7'h0,_GEN_1164};
  assign _T_25298 = {7'h0,_GEN_1165};
  assign _T_25300 = {7'h0,_GEN_1166};
  assign _T_25302 = {7'h0,_GEN_1167};
  assign _T_25304 = {7'h0,_GEN_1168};
  assign _T_25306 = {7'h0,_GEN_1169};
  assign _T_25308 = {7'h0,_GEN_1170};
  assign _T_25310 = {7'h0,_GEN_1171};
  assign _T_25312 = {7'h0,_GEN_1172};
  assign _T_25314 = {7'h0,_GEN_1173};
  assign _T_25316 = {7'h0,_GEN_1174};
  assign _T_25318 = {7'h0,_GEN_1175};
  assign _T_25320 = {7'h0,_GEN_1176};
  assign _T_25322 = {7'h0,_GEN_1177};
  assign _T_25324 = {7'h0,_GEN_1178};
  assign _T_25326 = {7'h0,_GEN_1179};
  assign _T_25328 = {7'h0,_GEN_1180};
  assign _T_25330 = {7'h0,_GEN_1181};
  assign _T_25332 = {7'h0,_GEN_1182};
  assign _T_25334 = {7'h0,_GEN_1183};
  assign _T_25336 = {7'h0,_GEN_1184};
  assign _T_25338 = {7'h0,_GEN_1185};
  assign _T_25340 = {7'h0,_GEN_1186};
  assign _T_25342 = {7'h0,_GEN_1187};
  assign _T_25344 = {7'h0,_GEN_1188};
  assign _T_25346 = {7'h0,_GEN_1189};
  assign _T_25348 = {7'h0,_GEN_1190};
  assign _T_25350 = {7'h0,_GEN_1191};
  assign _T_25352 = {7'h0,_GEN_1192};
  assign _T_25354 = {7'h0,_GEN_1193};
  assign _T_25356 = {7'h0,_GEN_1194};
  assign _T_25358 = {7'h0,_GEN_1195};
  assign _T_25360 = {7'h0,_GEN_1196};
  assign _T_25362 = {7'h0,_GEN_1197};
  assign _T_25364 = {7'h0,_GEN_1198};
  assign _T_25366 = {7'h0,_GEN_1199};
  assign _T_25368 = {7'h0,_GEN_1200};
  assign _T_25370 = {7'h0,_GEN_1201};
  assign _T_25372 = {7'h0,_GEN_1202};
  assign _T_25374 = {7'h0,_GEN_1203};
  assign _T_25376 = {7'h0,_GEN_1204};
  assign _T_25378 = {7'h0,_GEN_1205};
  assign _T_25380 = {7'h0,_GEN_1206};
  assign _T_25382 = {7'h0,_GEN_1207};
  assign _T_25384 = {7'h0,_GEN_1208};
  assign _T_25386 = {7'h0,_GEN_1209};
  assign _T_25388 = {7'h0,_GEN_1210};
  assign _T_25390 = {7'h0,_GEN_1211};
  assign _T_25392 = {7'h0,_GEN_1212};
  assign _T_25394 = {7'h0,_GEN_1213};
  assign _T_25396 = {7'h0,_GEN_1214};
  assign _T_25398 = {7'h0,_GEN_1215};
  assign _T_25400 = {7'h0,_GEN_1216};
  assign _T_25402 = {7'h0,_GEN_1217};
  assign _T_25404 = {7'h0,_GEN_1218};
  assign _T_25406 = {7'h0,_GEN_1219};
  assign _T_25408 = {7'h0,_GEN_1220};
  assign _T_25410 = {7'h0,_GEN_1221};
  assign _T_25412 = {7'h0,_GEN_1222};
  assign _T_25414 = {7'h0,_GEN_1223};
  assign _T_25416 = {7'h0,_GEN_1224};
  assign _T_25418 = {7'h0,_GEN_1225};
  assign _T_25420 = {7'h0,_GEN_1226};
  assign _T_25422 = {7'h0,_GEN_1227};
  assign _T_25424 = {7'h0,_GEN_1228};
  assign _T_25426 = {7'h0,_GEN_1229};
  assign _T_25428 = {7'h0,_GEN_1230};
  assign _T_25430 = {7'h0,_GEN_1231};
  assign _T_25432 = {7'h0,_GEN_1232};
  assign _T_25434 = {7'h0,_GEN_1233};
  assign _T_25436 = {7'h0,_GEN_1234};
  assign _T_25438 = {7'h0,_GEN_1235};
  assign _T_25440 = {7'h0,_GEN_1236};
  assign _T_25442 = {7'h0,_GEN_1237};
  assign _T_25444 = {7'h0,_GEN_1238};
  assign _T_25446 = {7'h0,_GEN_1239};
  assign _T_25448 = {7'h0,_GEN_1240};
  assign _T_25450 = {7'h0,_GEN_1241};
  assign _T_25452 = {7'h0,_GEN_1242};
  assign _T_25454 = {7'h0,_GEN_1243};
  assign _T_25456 = {7'h0,_GEN_1244};
  assign _T_25458 = {7'h0,_GEN_1245};
  assign _T_25460 = {7'h0,_GEN_1246};
  assign _T_25462 = {7'h0,_GEN_1247};
  assign _T_25464 = {7'h0,_GEN_1248};
  assign _T_25466 = {7'h0,_GEN_1249};
  assign _T_25468 = {7'h0,_GEN_1250};
  assign _T_25470 = {7'h0,_GEN_1251};
  assign _T_25472 = {7'h0,_GEN_1252};
  assign _T_25474 = {7'h0,_GEN_1253};
  assign _T_25476 = {7'h0,_GEN_1254};
  assign _T_25478 = {7'h0,_GEN_1255};
  assign _T_25480 = {7'h0,_GEN_1256};
  assign _T_25482 = {7'h0,_GEN_1257};
  assign _T_25484 = {7'h0,_GEN_1258};
  assign _T_25486 = {7'h0,_GEN_1259};
  assign _T_25488 = {7'h0,_GEN_1260};
  assign _T_25490 = {7'h0,_GEN_1261};
  assign _T_25492 = {7'h0,_GEN_1262};
  assign _T_25494 = {7'h0,_GEN_1263};
  assign _T_25496 = {7'h0,_GEN_1264};
  assign _T_25498 = {7'h0,_GEN_1265};
  assign _T_25500 = {7'h0,_GEN_1266};
  assign _T_25502 = {7'h0,_GEN_1267};
  assign _T_25504 = {7'h0,_GEN_1268};
  assign _T_25506 = {7'h0,_GEN_1269};
  assign _T_25508 = {7'h0,_GEN_1270};
  assign _T_25510 = {7'h0,_GEN_1271};
  assign _T_25512 = {7'h0,_GEN_1272};
  assign _T_25514 = {7'h0,_GEN_1273};
  assign _T_25516 = {7'h0,_GEN_1274};
  assign _T_25518 = {7'h0,_GEN_1275};
  assign _T_25520 = {7'h0,_GEN_1276};
  assign _T_25522 = {7'h0,_GEN_1277};
  assign _T_25524 = {7'h0,_GEN_1278};
  assign _T_25526 = {7'h0,_GEN_1279};
  assign _T_25528 = {7'h0,_GEN_1280};
  assign _T_25530 = {7'h0,_GEN_1281};
  assign _T_25532 = {7'h0,_GEN_1282};
  assign _T_25534 = {7'h0,_GEN_1283};
  assign _T_25536 = {7'h0,_GEN_1284};
  assign _T_25538 = {7'h0,_GEN_1285};
  assign _T_25540 = {7'h0,_GEN_1286};
  assign _T_25542 = {7'h0,_GEN_1287};
  assign _T_25544 = {7'h0,_GEN_1288};
  assign _T_25546 = {7'h0,_GEN_1289};
  assign _T_25548 = {7'h0,_GEN_1290};
  assign _T_25550 = {7'h0,_GEN_1291};
  assign _T_25552 = {7'h0,_GEN_1292};
  assign _T_25554 = {7'h0,_GEN_1293};
  assign _T_25556 = {7'h0,_GEN_1294};
  assign _T_25558 = {7'h0,_GEN_1295};
  assign _T_25560 = {7'h0,_GEN_1296};
  assign _T_25562 = {7'h0,_GEN_1297};
  assign _T_25564 = {7'h0,_GEN_1298};
  assign _T_25566 = {7'h0,_GEN_1299};
  assign _T_25568 = {7'h0,_GEN_1300};
  assign _T_25570 = {7'h0,_GEN_1301};
  assign _T_25572 = {7'h0,_GEN_1302};
  assign _T_25574 = {7'h0,_GEN_1303};
  assign _T_25576 = {7'h0,_GEN_1304};
  assign _T_25578 = {7'h0,_GEN_1305};
  assign _T_25580 = {7'h0,_GEN_1306};
  assign _T_25582 = {7'h0,_GEN_1307};
  assign _T_25584 = {7'h0,_GEN_1308};
  assign _T_25586 = {7'h0,_GEN_1309};
  assign _T_25588 = {7'h0,_GEN_1310};
  assign _T_25590 = {7'h0,_GEN_1311};
  assign _T_25592 = {7'h0,_GEN_1312};
  assign _T_25594 = {7'h0,_GEN_1313};
  assign _T_25596 = {7'h0,_GEN_1314};
  assign _T_25598 = {7'h0,_GEN_1315};
  assign _T_25600 = {7'h0,_GEN_1316};
  assign _T_25602 = {7'h0,_GEN_1317};
  assign _T_25604 = {7'h0,_GEN_1318};
  assign _T_25606 = {7'h0,_GEN_1319};
  assign _T_25608 = {7'h0,_GEN_1320};
  assign _T_25610 = {7'h0,_GEN_1321};
  assign _T_25612 = {7'h0,_GEN_1322};
  assign _T_25614 = {7'h0,_GEN_1323};
  assign _T_25616 = {7'h0,_GEN_1324};
  assign _T_25618 = {7'h0,_GEN_1325};
  assign _T_25620 = {7'h0,_GEN_1326};
  assign _T_25622 = {7'h0,_GEN_1327};
  assign _T_25624 = {7'h0,_GEN_1328};
  assign _T_25626 = {7'h0,_GEN_1329};
  assign _T_25628 = {7'h0,_GEN_1330};
  assign _T_25630 = {7'h0,_GEN_1331};
  assign _T_25632 = {7'h0,_GEN_1332};
  assign _T_25634 = {7'h0,_GEN_1333};
  assign _T_25636 = {7'h0,_GEN_1334};
  assign _T_25638 = {7'h0,_GEN_1335};
  assign _T_25640 = {7'h0,_GEN_1336};
  assign _T_25642 = {7'h0,_GEN_1337};
  assign _T_25644 = {7'h0,_GEN_1338};
  assign _T_25646 = {7'h0,_GEN_1339};
  assign _T_25648 = {7'h0,_GEN_1340};
  assign _T_25650 = {7'h0,_GEN_1341};
  assign _T_25652 = {7'h0,_GEN_1342};
  assign _T_25654 = {7'h0,_GEN_1343};
  assign _T_25656 = {7'h0,_GEN_1344};
  assign _T_25658 = {7'h0,_GEN_1345};
  assign _T_25660 = {7'h0,_GEN_1346};
  assign _T_25662 = {7'h0,_GEN_1347};
  assign _T_25664 = {7'h0,_GEN_1348};
  assign _T_25666 = {7'h0,_GEN_1349};
  assign _T_25668 = {7'h0,_GEN_1350};
  assign _T_25670 = {7'h0,_GEN_1351};
  assign _T_25672 = {7'h0,_GEN_1352};
  assign _T_25674 = {7'h0,_GEN_1353};
  assign _T_25676 = {7'h0,_GEN_1354};
  assign _T_25678 = {7'h0,_GEN_1355};
  assign _T_25680 = {7'h0,_GEN_1356};
  assign _T_25682 = {7'h0,_GEN_1357};
  assign _T_25684 = {7'h0,_GEN_1358};
  assign _T_25686 = {7'h0,_GEN_1359};
  assign _T_25688 = {7'h0,_GEN_1360};
  assign _T_25690 = {7'h0,_GEN_1361};
  assign _T_25692 = {7'h0,_GEN_1362};
  assign _T_25694 = {7'h0,_GEN_1363};
  assign _T_25696 = {7'h0,_GEN_1364};
  assign _T_25698 = {7'h0,_GEN_1365};
  assign _T_25700 = {7'h0,_GEN_1366};
  assign _T_25702 = {7'h0,_GEN_1367};
  assign _T_25704 = {7'h0,_GEN_1368};
  assign _T_25706 = {7'h0,_GEN_1369};
  assign _T_25708 = {7'h0,_GEN_1370};
  assign _T_25710 = {7'h0,_GEN_1371};
  assign _T_25712 = {7'h0,_GEN_1372};
  assign _T_25714 = {7'h0,_GEN_1373};
  assign _T_25716 = {7'h0,_GEN_1374};
  assign _T_25718 = {7'h0,_GEN_1375};
  assign _T_25720 = {7'h0,_GEN_1376};
  assign _T_25722 = {7'h0,_GEN_1377};
  assign _T_25724 = {7'h0,_GEN_1378};
  assign _T_25726 = {7'h0,_GEN_1379};
  assign _T_25728 = {7'h0,_GEN_1380};
  assign _T_25730 = {7'h0,_GEN_1381};
  assign _T_25732 = {7'h0,_GEN_1382};
  assign _T_25734 = {7'h0,_GEN_1383};
  assign _T_25736 = {7'h0,_GEN_1384};
  assign _T_25738 = {7'h0,_GEN_1385};
  assign _T_25740 = {7'h0,_GEN_1386};
  assign _T_25742 = {7'h0,_GEN_1387};
  assign _T_25744 = {7'h0,_GEN_1388};
  assign _T_25746 = {7'h0,_GEN_1389};
  assign _T_25748 = {7'h0,_GEN_1390};
  assign _T_25750 = {7'h0,_GEN_1391};
  assign _T_25752 = {7'h0,_GEN_1392};
  assign _T_25754 = {7'h0,_GEN_1393};
  assign _T_25756 = {7'h0,_GEN_1394};
  assign _T_25758 = {7'h0,_GEN_1395};
  assign _T_25760 = {7'h0,_GEN_1396};
  assign _T_25762 = {7'h0,_GEN_1397};
  assign _T_25764 = {7'h0,_GEN_1398};
  assign _T_25766 = {7'h0,_GEN_1399};
  assign _T_25768 = {7'h0,_GEN_1400};
  assign _T_25770 = {7'h0,_GEN_1401};
  assign _T_25772 = {7'h0,_GEN_1402};
  assign _T_25774 = {7'h0,_GEN_1403};
  assign _T_25776 = {7'h0,_GEN_1404};
  assign _T_25778 = {7'h0,_GEN_1405};
  assign _T_25780 = {7'h0,_GEN_1406};
  assign _T_25782 = {7'h0,_GEN_1407};
  assign _T_25784 = {7'h0,_GEN_1408};
  assign _T_25786 = {7'h0,_GEN_1409};
  assign _T_25788 = {7'h0,_GEN_1410};
  assign _T_25790 = {7'h0,_GEN_1411};
  assign _T_25792 = {7'h0,_GEN_1412};
  assign _T_25899 = io_hart_in_0_a_bits_opcode == 3'h4;
  assign _T_25900 = io_hart_in_0_a_bits_address[11:2];
  assign _T_25901 = {io_hart_in_0_a_bits_source,io_hart_in_0_a_bits_size};
  assign _T_26947 = _T_25900 ^ 10'h16d;
  assign _T_26948 = _T_26947 & 10'h200;
  assign _T_26950 = _T_26948 == 10'h0;
  assign _T_26956 = _T_25900 ^ 10'h1df;
  assign _T_26957 = _T_26956 & 10'h200;
  assign _T_26959 = _T_26957 == 10'h0;
  assign _T_26965 = _T_25900 ^ 10'h15b;
  assign _T_26966 = _T_26965 & 10'h200;
  assign _T_26968 = _T_26966 == 10'h0;
  assign _T_26974 = _T_25900 ^ 10'h14d;
  assign _T_26975 = _T_26974 & 10'h200;
  assign _T_26977 = _T_26975 == 10'h0;
  assign _T_26983 = _T_25900 ^ 10'h206;
  assign _T_26984 = _T_26983 & 10'h200;
  assign _T_26986 = _T_26984 == 10'h0;
  assign _T_26992 = _T_25900 ^ 10'h1d4;
  assign _T_26993 = _T_26992 & 10'h200;
  assign _T_26995 = _T_26993 == 10'h0;
  assign _T_27001 = _T_25900 ^ 10'h1e1;
  assign _T_27002 = _T_27001 & 10'h200;
  assign _T_27004 = _T_27002 == 10'h0;
  assign _T_27010 = _T_25900 ^ 10'h160;
  assign _T_27011 = _T_27010 & 10'h200;
  assign _T_27013 = _T_27011 == 10'h0;
  assign _T_27019 = _T_25900 ^ 10'h198;
  assign _T_27020 = _T_27019 & 10'h200;
  assign _T_27022 = _T_27020 == 10'h0;
  assign _T_27028 = _T_25900 ^ 10'h20b;
  assign _T_27029 = _T_27028 & 10'h200;
  assign _T_27031 = _T_27029 == 10'h0;
  assign _T_27037 = _T_25900 ^ 10'hd9;
  assign _T_27038 = _T_27037 & 10'h200;
  assign _T_27040 = _T_27038 == 10'h0;
  assign _T_27046 = _T_25900 ^ 10'h114;
  assign _T_27047 = _T_27046 & 10'h200;
  assign _T_27049 = _T_27047 == 10'h0;
  assign _T_27055 = _T_25900 ^ 10'h134;
  assign _T_27056 = _T_27055 & 10'h200;
  assign _T_27058 = _T_27056 == 10'h0;
  assign _T_27064 = _T_25900 ^ 10'h1c1;
  assign _T_27065 = _T_27064 & 10'h200;
  assign _T_27067 = _T_27065 == 10'h0;
  assign _T_27073 = _T_25900 ^ 10'h17b;
  assign _T_27074 = _T_27073 & 10'h200;
  assign _T_27076 = _T_27074 == 10'h0;
  assign _T_27082 = _T_25900 ^ 10'h1b8;
  assign _T_27083 = _T_27082 & 10'h200;
  assign _T_27085 = _T_27083 == 10'h0;
  assign _T_27091 = _T_25900 ^ 10'h1ff;
  assign _T_27092 = _T_27091 & 10'h200;
  assign _T_27094 = _T_27092 == 10'h0;
  assign _T_27100 = _T_25900 ^ 10'h10d;
  assign _T_27101 = _T_27100 & 10'h200;
  assign _T_27103 = _T_27101 == 10'h0;
  assign _T_27109 = _T_25900 ^ 10'h181;
  assign _T_27110 = _T_27109 & 10'h200;
  assign _T_27112 = _T_27110 == 10'h0;
  assign _T_27118 = _T_25900 ^ 10'h180;
  assign _T_27119 = _T_27118 & 10'h200;
  assign _T_27121 = _T_27119 == 10'h0;
  assign _T_27127 = _T_25900 ^ 10'h215;
  assign _T_27128 = _T_27127 & 10'h200;
  assign _T_27130 = _T_27128 == 10'h0;
  assign _T_27136 = _T_25900 ^ 10'h1f4;
  assign _T_27137 = _T_27136 & 10'h200;
  assign _T_27139 = _T_27137 == 10'h0;
  assign _T_27145 = _T_25900 ^ 10'h1d8;
  assign _T_27146 = _T_27145 & 10'h200;
  assign _T_27148 = _T_27146 == 10'h0;
  assign _T_27154 = _T_25900 ^ 10'h154;
  assign _T_27155 = _T_27154 & 10'h200;
  assign _T_27157 = _T_27155 == 10'h0;
  assign _T_27163 = _T_25900 ^ 10'h194;
  assign _T_27164 = _T_27163 & 10'h200;
  assign _T_27166 = _T_27164 == 10'h0;
  assign _T_27172 = _T_25900 ^ 10'h1a1;
  assign _T_27173 = _T_27172 & 10'h200;
  assign _T_27175 = _T_27173 == 10'h0;
  assign _T_27181 = _T_25900 ^ 10'h120;
  assign _T_27182 = _T_27181 & 10'h200;
  assign _T_27184 = _T_27182 == 10'h0;
  assign _T_27190 = _T_25900 ^ 10'h12d;
  assign _T_27191 = _T_27190 & 10'h200;
  assign _T_27193 = _T_27191 == 10'h0;
  assign _T_27199 = _T_25900 ^ 10'h140;
  assign _T_27200 = _T_27199 & 10'h200;
  assign _T_27202 = _T_27200 == 10'h0;
  assign _T_27208 = _T_25900 ^ 10'h1b4;
  assign _T_27209 = _T_27208 & 10'h200;
  assign _T_27211 = _T_27209 == 10'h0;
  assign _T_27217 = _T_25900 ^ 10'h101;
  assign _T_27218 = _T_27217 & 10'h200;
  assign _T_27220 = _T_27218 == 10'h0;
  assign _T_27226 = _T_25900 ^ 10'h185;
  assign _T_27227 = _T_27226 & 10'h200;
  assign _T_27229 = _T_27227 == 10'h0;
  assign _T_27235 = _T_25900 ^ 10'h174;
  assign _T_27236 = _T_27235 & 10'h200;
  assign _T_27238 = _T_27236 == 10'h0;
  assign _T_27244 = _T_25900 ^ 10'h1f8;
  assign _T_27245 = _T_27244 & 10'h200;
  assign _T_27247 = _T_27245 == 10'h0;
  assign _T_27253 = _T_25900 ^ 10'h158;
  assign _T_27254 = _T_27253 & 10'h200;
  assign _T_27256 = _T_27254 == 10'h0;
  assign _T_27262 = _T_25900 ^ 10'h165;
  assign _T_27263 = _T_27262 & 10'h200;
  assign _T_27265 = _T_27263 == 10'h0;
  assign _T_27271 = _T_25900 ^ 10'h1cc;
  assign _T_27272 = _T_27271 & 10'h200;
  assign _T_27274 = _T_27272 == 10'h0;
  assign _T_27280 = _T_25900 ^ 10'h1a5;
  assign _T_27281 = _T_27280 & 10'h200;
  assign _T_27283 = _T_27281 == 10'h0;
  assign _T_27289 = _T_25900 ^ 10'h11c;
  assign _T_27290 = _T_27289 & 10'h200;
  assign _T_27292 = _T_27290 == 10'h0;
  assign _T_27298 = _T_25900 ^ 10'h1a0;
  assign _T_27299 = _T_27298 & 10'h200;
  assign _T_27301 = _T_27299 == 10'h0;
  assign _T_27307 = _T_25900 ^ 10'h145;
  assign _T_27308 = _T_27307 & 10'h200;
  assign _T_27310 = _T_27308 == 10'h0;
  assign _T_27316 = _T_25900 ^ 10'h121;
  assign _T_27317 = _T_27316 & 10'h200;
  assign _T_27319 = _T_27317 == 10'h0;
  assign _T_27325 = _T_25900 ^ 10'h1c0;
  assign _T_27326 = _T_27325 & 10'h200;
  assign _T_27328 = _T_27326 == 10'h0;
  assign _T_27334 = _T_25900 ^ 10'h13c;
  assign _T_27335 = _T_27334 & 10'h200;
  assign _T_27337 = _T_27335 == 10'h0;
  assign _T_27343 = _T_25900 ^ 10'h105;
  assign _T_27344 = _T_27343 & 10'h200;
  assign _T_27346 = _T_27344 == 10'h0;
  assign _T_27352 = _T_25900 ^ 10'hd8;
  assign _T_27353 = _T_27352 & 10'h200;
  assign _T_27355 = _T_27353 == 10'h0;
  assign _T_27361 = _T_25900 ^ 10'h1db;
  assign _T_27362 = _T_27361 & 10'h200;
  assign _T_27364 = _T_27362 == 10'h0;
  assign _T_27370 = _T_25900 ^ 10'h1ec;
  assign _T_27371 = _T_27370 & 10'h200;
  assign _T_27373 = _T_27371 == 10'h0;
  assign _T_27379 = _T_25900 ^ 10'h1bb;
  assign _T_27380 = _T_27379 & 10'h200;
  assign _T_27382 = _T_27380 == 10'h0;
  assign _T_27388 = _T_25900 ^ 10'h141;
  assign _T_27389 = _T_27388 & 10'h200;
  assign _T_27391 = _T_27389 == 10'h0;
  assign _T_27397 = _T_25900 ^ 10'h178;
  assign _T_27398 = _T_27397 & 10'h200;
  assign _T_27400 = _T_27398 == 10'h0;
  assign _T_27406 = _T_25900 ^ 10'hd3;
  assign _T_27407 = _T_27406 & 10'h200;
  assign _T_27409 = _T_27407 == 10'h0;
  assign _T_27415 = _T_25900 ^ 10'h1e5;
  assign _T_27416 = _T_27415 & 10'h200;
  assign _T_27418 = _T_27416 == 10'h0;
  assign _T_27424 = _T_25900 ^ 10'h202;
  assign _T_27425 = _T_27424 & 10'h200;
  assign _T_27427 = _T_27425 == 10'h0;
  assign _T_27433 = _T_25900 ^ 10'h15c;
  assign _T_27434 = _T_27433 & 10'h200;
  assign _T_27436 = _T_27434 == 10'h0;
  assign _T_27442 = _T_25900 ^ 10'h161;
  assign _T_27443 = _T_27442 & 10'h200;
  assign _T_27445 = _T_27443 == 10'h0;
  assign _T_27451 = _T_25900 ^ 10'h1e0;
  assign _T_27452 = _T_27451 & 10'h200;
  assign _T_27454 = _T_27452 == 10'h0;
  assign _T_27460 = _T_25900 ^ 10'h18d;
  assign _T_27461 = _T_27460 & 10'h200;
  assign _T_27463 = _T_27461 == 10'h0;
  assign _T_27469 = _T_25900 ^ 10'h118;
  assign _T_27470 = _T_27469 & 10'h200;
  assign _T_27472 = _T_27470 == 10'h0;
  assign _T_27478 = _T_25900 ^ 10'hdd;
  assign _T_27479 = _T_27478 & 10'h200;
  assign _T_27481 = _T_27479 == 10'h0;
  assign _T_27487 = _T_25900 ^ 10'h125;
  assign _T_27488 = _T_27487 & 10'h200;
  assign _T_27490 = _T_27488 == 10'h0;
  assign _T_27496 = _T_25900 ^ 10'h1c5;
  assign _T_27497 = _T_27496 & 10'h200;
  assign _T_27499 = _T_27497 == 10'h0;
  assign _T_27505 = _T_25900 ^ 10'h18c;
  assign _T_27506 = _T_27505 & 10'h200;
  assign _T_27508 = _T_27506 == 10'h0;
  assign _T_27514 = _T_25900 ^ 10'h19b;
  assign _T_27515 = _T_27514 & 10'h200;
  assign _T_27517 = _T_27515 == 10'h0;
  assign _T_27523 = _T_25900 ^ 10'h1ac;
  assign _T_27524 = _T_27523 & 10'h200;
  assign _T_27526 = _T_27524 == 10'h0;
  assign _T_27532 = _T_25900 ^ 10'h109;
  assign _T_27533 = _T_27532 & 10'h200;
  assign _T_27535 = _T_27533 == 10'h0;
  assign _T_27541 = _T_25900 ^ 10'h1fb;
  assign _T_27542 = _T_27541 & 10'h200;
  assign _T_27544 = _T_27542 == 10'h0;
  assign _T_27550 = _T_25900 ^ 10'h20f;
  assign _T_27551 = _T_27550 & 10'h200;
  assign _T_27553 = _T_27551 == 10'h0;
  assign _T_27559 = _T_25900 ^ 10'h138;
  assign _T_27560 = _T_27559 & 10'h200;
  assign _T_27562 = _T_27560 == 10'h0;
  assign _T_27568 = _T_25900 ^ 10'hce;
  assign _T_27569 = _T_27568 & 10'h200;
  assign _T_27571 = _T_27569 == 10'h0;
  assign _T_27577 = _T_25900 ^ 10'h133;
  assign _T_27578 = _T_27577 & 10'h200;
  assign _T_27580 = _T_27578 == 10'h0;
  assign _T_27586 = _T_25900 ^ 10'h124;
  assign _T_27587 = _T_27586 & 10'h200;
  assign _T_27589 = _T_27587 == 10'h0;
  assign _T_27595 = _T_25900 ^ 10'h1c4;
  assign _T_27596 = _T_27595 & 10'h200;
  assign _T_27598 = _T_27596 == 10'h0;
  assign _T_27604 = _T_25900 ^ 10'h17c;
  assign _T_27605 = _T_27604 & 10'h200;
  assign _T_27607 = _T_27605 == 10'h0;
  assign _T_27613 = _T_25900 ^ 10'h200;
  assign _T_27614 = _T_27613 & 10'h200;
  assign _T_27616 = _T_27614 == 10'h0;
  assign _T_27622 = _T_25900 ^ 10'h1b7;
  assign _T_27623 = _T_27622 & 10'h200;
  assign _T_27625 = _T_27623 == 10'h0;
  assign _T_27631 = _T_25900 ^ 10'h10e;
  assign _T_27632 = _T_27631 & 10'h200;
  assign _T_27634 = _T_27632 == 10'h0;
  assign _T_27640 = _T_25900 ^ 10'h211;
  assign _T_27641 = _T_27640 & 10'h200;
  assign _T_27643 = _T_27641 == 10'h0;
  assign _T_27649 = _T_25900 ^ 10'h17d;
  assign _T_27650 = _T_27649 & 10'h200;
  assign _T_27652 = _T_27650 == 10'h0;
  assign _T_27658 = _T_25900 ^ 10'hdc;
  assign _T_27659 = _T_27658 & 10'h200;
  assign _T_27661 = _T_27659 == 10'h0;
  assign _T_27667 = _T_25900 ^ 10'h16e;
  assign _T_27668 = _T_27667 & 10'h200;
  assign _T_27670 = _T_27668 == 10'h0;
  assign _T_27676 = _T_25900 ^ 10'h216;
  assign _T_27677 = _T_27676 & 10'h200;
  assign _T_27679 = _T_27677 == 10'h0;
  assign _T_27685 = _T_25900 ^ 10'h14e;
  assign _T_27686 = _T_27685 & 10'h200;
  assign _T_27688 = _T_27686 == 10'h0;
  assign _T_27694 = _T_25900 ^ 10'h12e;
  assign _T_27695 = _T_27694 & 10'h200;
  assign _T_27697 = _T_27695 == 10'h0;
  assign _T_27703 = _T_25900 ^ 10'h104;
  assign _T_27704 = _T_27703 & 10'h200;
  assign _T_27706 = _T_27704 == 10'h0;
  assign _T_27712 = _T_25900 ^ 10'h15d;
  assign _T_27713 = _T_27712 & 10'h200;
  assign _T_27715 = _T_27713 == 10'h0;
  assign _T_27721 = _T_25900 ^ 10'h188;
  assign _T_27722 = _T_27721 & 10'h200;
  assign _T_27724 = _T_27722 == 10'h0;
  assign _T_27730 = _T_25900 ^ 10'h129;
  assign _T_27731 = _T_27730 & 10'h200;
  assign _T_27733 = _T_27731 == 10'h0;
  assign _T_27739 = _T_25900 ^ 10'h1a8;
  assign _T_27740 = _T_27739 & 10'h200;
  assign _T_27742 = _T_27740 == 10'h0;
  assign _T_27748 = _T_25900 ^ 10'hc0;
  assign _T_27749 = _T_27748 & 10'h200;
  assign _T_27751 = _T_27749 == 10'h0;
  assign _T_27757 = _T_25900 ^ 10'h197;
  assign _T_27758 = _T_27757 & 10'h200;
  assign _T_27760 = _T_27758 == 10'h0;
  assign _T_27766 = _T_25900 ^ 10'h1ad;
  assign _T_27767 = _T_27766 & 10'h200;
  assign _T_27769 = _T_27767 == 10'h0;
  assign _T_27775 = _T_25900 ^ 10'h113;
  assign _T_27776 = _T_27775 & 10'h200;
  assign _T_27778 = _T_27776 == 10'h0;
  assign _T_27784 = _T_25900 ^ 10'h1d3;
  assign _T_27785 = _T_27784 & 10'h200;
  assign _T_27787 = _T_27785 == 10'h0;
  assign _T_27793 = _T_25900 ^ 10'h1e4;
  assign _T_27794 = _T_27793 & 10'h200;
  assign _T_27796 = _T_27794 == 10'h0;
  assign _T_27802 = _T_25900 ^ 10'h169;
  assign _T_27803 = _T_27802 & 10'h200;
  assign _T_27805 = _T_27803 == 10'h0;
  assign _T_27811 = _T_25900 ^ 10'h41;
  assign _T_27812 = _T_27811 & 10'h200;
  assign _T_27814 = _T_27812 == 10'h0;
  assign _T_27820 = _T_25900 ^ 10'h1b3;
  assign _T_27821 = _T_27820 & 10'h200;
  assign _T_27823 = _T_27821 == 10'h0;
  assign _T_27829 = _T_25900 ^ 10'h149;
  assign _T_27830 = _T_27829 & 10'h200;
  assign _T_27832 = _T_27830 == 10'h0;
  assign _T_27838 = _T_25900 ^ 10'h20a;
  assign _T_27839 = _T_27838 & 10'h200;
  assign _T_27841 = _T_27839 == 10'h0;
  assign _T_27847 = _T_25900 ^ 10'h1cd;
  assign _T_27848 = _T_27847 & 10'h200;
  assign _T_27850 = _T_27848 == 10'h0;
  assign _T_27856 = _T_25900 ^ 10'h1ed;
  assign _T_27857 = _T_27856 & 10'h200;
  assign _T_27859 = _T_27857 == 10'h0;
  assign _T_27865 = _T_25900 ^ 10'h1c8;
  assign _T_27866 = _T_27865 & 10'h200;
  assign _T_27868 = _T_27866 == 10'h0;
  assign _T_27874 = _T_25900 ^ 10'h144;
  assign _T_27875 = _T_27874 & 10'h200;
  assign _T_27877 = _T_27875 == 10'h0;
  assign _T_27883 = _T_25900 ^ 10'h11d;
  assign _T_27884 = _T_27883 & 10'h200;
  assign _T_27886 = _T_27884 == 10'h0;
  assign _T_27892 = _T_25900 ^ 10'he0;
  assign _T_27893 = _T_27892 & 10'h200;
  assign _T_27895 = _T_27893 == 10'h0;
  assign _T_27901 = _T_25900 ^ 10'h207;
  assign _T_27902 = _T_27901 & 10'h200;
  assign _T_27904 = _T_27902 == 10'h0;
  assign _T_27910 = _T_25900 ^ 10'h13d;
  assign _T_27911 = _T_27910 & 10'h200;
  assign _T_27913 = _T_27911 == 10'h0;
  assign _T_27919 = _T_25900 ^ 10'h193;
  assign _T_27920 = _T_27919 & 10'h200;
  assign _T_27922 = _T_27920 == 10'h0;
  assign _T_27928 = _T_25900 ^ 10'h184;
  assign _T_27929 = _T_27928 & 10'h200;
  assign _T_27931 = _T_27929 == 10'h0;
  assign _T_27937 = _T_25900 ^ 10'h164;
  assign _T_27938 = _T_27937 & 10'h200;
  assign _T_27940 = _T_27938 == 10'h0;
  assign _T_27946 = _T_25900 ^ 10'h1a4;
  assign _T_27947 = _T_27946 & 10'h200;
  assign _T_27949 = _T_27947 == 10'h0;
  assign _T_27955 = _T_25900 ^ 10'h1f3;
  assign _T_27956 = _T_27955 & 10'h200;
  assign _T_27958 = _T_27956 == 10'h0;
  assign _T_27964 = _T_25900 ^ 10'h148;
  assign _T_27965 = _T_27964 & 10'h200;
  assign _T_27967 = _T_27965 == 10'h0;
  assign _T_27973 = _T_25900 ^ 10'h1d7;
  assign _T_27974 = _T_27973 & 10'h200;
  assign _T_27976 = _T_27974 == 10'h0;
  assign _T_27982 = _T_25900 ^ 10'h100;
  assign _T_27983 = _T_27982 & 10'h200;
  assign _T_27985 = _T_27983 == 10'h0;
  assign _T_27991 = _T_25900 ^ 10'h1e8;
  assign _T_27992 = _T_27991 & 10'h200;
  assign _T_27994 = _T_27992 == 10'h0;
  assign _T_28000 = _T_25900 ^ 10'h153;
  assign _T_28001 = _T_28000 & 10'h200;
  assign _T_28003 = _T_28001 == 10'h0;
  assign _T_28009 = _T_25900 ^ 10'h1dc;
  assign _T_28010 = _T_28009 & 10'h200;
  assign _T_28012 = _T_28010 == 10'h0;
  assign _T_28018 = _T_25900 ^ 10'h20e;
  assign _T_28019 = _T_28018 & 10'h200;
  assign _T_28021 = _T_28019 == 10'h0;
  assign _T_28027 = _T_25900 ^ 10'h1e9;
  assign _T_28028 = _T_28027 & 10'h200;
  assign _T_28030 = _T_28028 == 10'h0;
  assign _T_28036 = _T_25900 ^ 10'hd4;
  assign _T_28037 = _T_28036 & 10'h200;
  assign _T_28039 = _T_28037 == 10'h0;
  assign _T_28045 = _T_25900 ^ 10'h189;
  assign _T_28046 = _T_28045 & 10'h200;
  assign _T_28048 = _T_28046 == 10'h0;
  assign _T_28054 = _T_25900 ^ 10'h203;
  assign _T_28055 = _T_28054 & 10'h200;
  assign _T_28057 = _T_28055 == 10'h0;
  assign _T_28063 = _T_25900 ^ 10'h1c9;
  assign _T_28064 = _T_28063 & 10'h200;
  assign _T_28066 = _T_28064 == 10'h0;
  assign _T_28072 = _T_25900 ^ 10'h173;
  assign _T_28073 = _T_28072 & 10'h200;
  assign _T_28075 = _T_28073 == 10'h0;
  assign _T_28081 = _T_25900 ^ 10'h1f7;
  assign _T_28082 = _T_28081 & 10'h200;
  assign _T_28084 = _T_28082 == 10'h0;
  assign _T_28090 = _T_25900 ^ 10'h157;
  assign _T_28091 = _T_28090 & 10'h200;
  assign _T_28093 = _T_28091 == 10'h0;
  assign _T_28099 = _T_25900 ^ 10'h10a;
  assign _T_28100 = _T_28099 & 10'h200;
  assign _T_28102 = _T_28100 == 10'h0;
  assign _T_28108 = _T_25900 ^ 10'h168;
  assign _T_28109 = _T_28108 & 10'h200;
  assign _T_28111 = _T_28109 == 10'h0;
  assign _T_28117 = _T_25900 ^ 10'h1fc;
  assign _T_28118 = _T_28117 & 10'h200;
  assign _T_28120 = _T_28118 == 10'h0;
  assign _T_28126 = _T_25900 ^ 10'h137;
  assign _T_28127 = _T_28126 & 10'h200;
  assign _T_28129 = _T_28127 == 10'h0;
  assign _T_28135 = _T_25900 ^ 10'h18e;
  assign _T_28136 = _T_28135 & 10'h200;
  assign _T_28138 = _T_28136 == 10'h0;
  assign _T_28144 = _T_25900 ^ 10'h212;
  assign _T_28145 = _T_28144 & 10'h200;
  assign _T_28147 = _T_28145 == 10'h0;
  assign _T_28153 = _T_25900 ^ 10'h12a;
  assign _T_28154 = _T_28153 & 10'h200;
  assign _T_28156 = _T_28154 == 10'h0;
  assign _T_28162 = _T_25900 ^ 10'h19c;
  assign _T_28163 = _T_28162 & 10'h200;
  assign _T_28165 = _T_28163 == 10'h0;
  assign _T_28171 = _T_25900 ^ 10'h1a9;
  assign _T_28172 = _T_28171 & 10'h200;
  assign _T_28174 = _T_28172 == 10'h0;
  assign _T_28180 = _T_25900 ^ 10'h201;
  assign _T_28181 = _T_28180 & 10'h200;
  assign _T_28183 = _T_28181 == 10'h0;
  assign _T_28189 = _T_25900 ^ 10'h1ae;
  assign _T_28190 = _T_28189 & 10'h200;
  assign _T_28192 = _T_28190 == 10'h0;
  assign _T_28198 = _T_25900 ^ 10'h108;
  assign _T_28199 = _T_28198 & 10'h200;
  assign _T_28201 = _T_28199 == 10'h0;
  assign _T_28207 = _T_25900 ^ 10'h117;
  assign _T_28208 = _T_28207 & 10'h200;
  assign _T_28210 = _T_28208 == 10'h0;
  assign _T_28216 = _T_25900 ^ 10'h40;
  assign _T_28217 = _T_28216 & 10'h200;
  assign _T_28219 = _T_28217 == 10'h0;
  assign _T_28225 = _T_25900 ^ 10'h128;
  assign _T_28226 = _T_28225 & 10'h200;
  assign _T_28228 = _T_28226 == 10'h0;
  assign _T_28234 = _T_25900 ^ 10'h1bc;
  assign _T_28235 = _T_28234 & 10'h200;
  assign _T_28237 = _T_28235 == 10'h0;
  assign _T_28243 = _T_25900 ^ 10'h177;
  assign _T_28244 = _T_28243 & 10'h200;
  assign _T_28246 = _T_28244 == 10'h0;
  assign _T_28252 = _T_25900 ^ 10'h1a7;
  assign _T_28253 = _T_28252 & 10'h200;
  assign _T_28255 = _T_28253 == 10'h0;
  assign _T_28261 = _T_25900 ^ 10'h192;
  assign _T_28262 = _T_28261 & 10'h200;
  assign _T_28264 = _T_28262 == 10'h0;
  assign _T_28270 = _T_25900 ^ 10'h11e;
  assign _T_28271 = _T_28270 & 10'h200;
  assign _T_28273 = _T_28271 == 10'h0;
  assign _T_28279 = _T_25900 ^ 10'h123;
  assign _T_28280 = _T_28279 & 10'h200;
  assign _T_28282 = _T_28280 == 10'h0;
  assign _T_28288 = _T_25900 ^ 10'h119;
  assign _T_28289 = _T_28288 & 10'h200;
  assign _T_28291 = _T_28289 == 10'h0;
  assign _T_28297 = _T_25900 ^ 10'h103;
  assign _T_28298 = _T_28297 & 10'h200;
  assign _T_28300 = _T_28298 == 10'h0;
  assign _T_28306 = _T_25900 ^ 10'h19d;
  assign _T_28307 = _T_28306 & 10'h200;
  assign _T_28309 = _T_28307 == 10'h0;
  assign _T_28315 = _T_25900 ^ 10'h187;
  assign _T_28316 = _T_28315 & 10'h200;
  assign _T_28318 = _T_28316 == 10'h0;
  assign _T_28324 = _T_25900 ^ 10'h1bd;
  assign _T_28325 = _T_28324 & 10'h200;
  assign _T_28327 = _T_28325 == 10'h0;
  assign _T_28333 = _T_25900 ^ 10'h17e;
  assign _T_28334 = _T_28333 & 10'h200;
  assign _T_28336 = _T_28334 == 10'h0;
  assign _T_28342 = _T_25900 ^ 10'h139;
  assign _T_28343 = _T_28342 & 10'h200;
  assign _T_28345 = _T_28343 == 10'h0;
  assign _T_28351 = _T_25900 ^ 10'h1f2;
  assign _T_28352 = _T_28351 & 10'h200;
  assign _T_28354 = _T_28352 == 10'h0;
  assign _T_28360 = _T_25900 ^ 10'h1d2;
  assign _T_28361 = _T_28360 & 10'h200;
  assign _T_28363 = _T_28361 == 10'h0;
  assign _T_28369 = _T_25900 ^ 10'h14f;
  assign _T_28370 = _T_28369 & 10'h200;
  assign _T_28372 = _T_28370 == 10'h0;
  assign _T_28378 = _T_25900 ^ 10'h15e;
  assign _T_28379 = _T_28378 & 10'h200;
  assign _T_28381 = _T_28379 == 10'h0;
  assign _T_28387 = _T_25900 ^ 10'h196;
  assign _T_28388 = _T_28387 & 10'h200;
  assign _T_28390 = _T_28388 == 10'h0;
  assign _T_28396 = _T_25900 ^ 10'hdb;
  assign _T_28397 = _T_28396 & 10'h200;
  assign _T_28399 = _T_28397 == 10'h0;
  assign _T_28405 = _T_25900 ^ 10'h112;
  assign _T_28406 = _T_28405 & 10'h200;
  assign _T_28408 = _T_28406 == 10'h0;
  assign _T_28414 = _T_25900 ^ 10'h1a3;
  assign _T_28415 = _T_28414 & 10'h200;
  assign _T_28417 = _T_28415 == 10'h0;
  assign _T_28423 = _T_25900 ^ 10'h179;
  assign _T_28424 = _T_28423 & 10'h200;
  assign _T_28426 = _T_28424 == 10'h0;
  assign _T_28432 = _T_25900 ^ 10'h16a;
  assign _T_28433 = _T_28432 & 10'h200;
  assign _T_28435 = _T_28433 == 10'h0;
  assign _T_28441 = _T_25900 ^ 10'h1c3;
  assign _T_28442 = _T_28441 & 10'h200;
  assign _T_28444 = _T_28442 == 10'h0;
  assign _T_28450 = _T_25900 ^ 10'h13e;
  assign _T_28451 = _T_28450 & 10'h200;
  assign _T_28453 = _T_28451 == 10'h0;
  assign _T_28459 = _T_25900 ^ 10'h1fd;
  assign _T_28460 = _T_28459 & 10'h200;
  assign _T_28462 = _T_28460 == 10'h0;
  assign _T_28468 = _T_25900 ^ 10'h1b2;
  assign _T_28469 = _T_28468 & 10'h200;
  assign _T_28471 = _T_28469 == 10'h0;
  assign _T_28477 = _T_25900 ^ 10'h12f;
  assign _T_28478 = _T_28477 & 10'h200;
  assign _T_28480 = _T_28478 == 10'h0;
  assign _T_28486 = _T_25900 ^ 10'h10f;
  assign _T_28487 = _T_28486 & 10'h200;
  assign _T_28489 = _T_28487 == 10'h0;
  assign _T_28495 = _T_25900 ^ 10'hd0;
  assign _T_28496 = _T_28495 & 10'h200;
  assign _T_28498 = _T_28496 == 10'h0;
  assign _T_28504 = _T_25900 ^ 10'h1dd;
  assign _T_28505 = _T_28504 & 10'h200;
  assign _T_28507 = _T_28505 == 10'h0;
  assign _T_28513 = _T_25900 ^ 10'h183;
  assign _T_28514 = _T_28513 & 10'h200;
  assign _T_28516 = _T_28514 == 10'h0;
  assign _T_28522 = _T_25900 ^ 10'h1ee;
  assign _T_28523 = _T_28522 & 10'h200;
  assign _T_28525 = _T_28523 == 10'h0;
  assign _T_28531 = _T_25900 ^ 10'h159;
  assign _T_28532 = _T_28531 & 10'h200;
  assign _T_28534 = _T_28532 == 10'h0;
  assign _T_28540 = _T_25900 ^ 10'h16f;
  assign _T_28541 = _T_28540 & 10'h200;
  assign _T_28543 = _T_28541 == 10'h0;
  assign _T_28549 = _T_25900 ^ 10'h217;
  assign _T_28550 = _T_28549 & 10'h200;
  assign _T_28552 = _T_28550 == 10'h0;
  assign _T_28558 = _T_25900 ^ 10'h143;
  assign _T_28559 = _T_28558 & 10'h200;
  assign _T_28561 = _T_28559 == 10'h0;
  assign _T_28567 = _T_25900 ^ 10'hd5;
  assign _T_28568 = _T_28567 & 10'h200;
  assign _T_28570 = _T_28568 == 10'h0;
  assign _T_28576 = _T_25900 ^ 10'h1e3;
  assign _T_28577 = _T_28576 & 10'h200;
  assign _T_28579 = _T_28577 == 10'h0;
  assign _T_28585 = _T_25900 ^ 10'h208;
  assign _T_28586 = _T_28585 & 10'h200;
  assign _T_28588 = _T_28586 == 10'h0;
  assign _T_28594 = _T_25900 ^ 10'h42;
  assign _T_28595 = _T_28594 & 10'h200;
  assign _T_28597 = _T_28595 == 10'h0;
  assign _T_28603 = _T_25900 ^ 10'h14a;
  assign _T_28604 = _T_28603 & 10'h200;
  assign _T_28606 = _T_28604 == 10'h0;
  assign _T_28612 = _T_25900 ^ 10'h1ce;
  assign _T_28613 = _T_28612 & 10'h200;
  assign _T_28615 = _T_28613 == 10'h0;
  assign _T_28621 = _T_25900 ^ 10'h209;
  assign _T_28622 = _T_28621 & 10'h200;
  assign _T_28624 = _T_28622 == 10'h0;
  assign _T_28630 = _T_25900 ^ 10'h18f;
  assign _T_28631 = _T_28630 & 10'h200;
  assign _T_28633 = _T_28631 == 10'h0;
  assign _T_28639 = _T_25900 ^ 10'h116;
  assign _T_28640 = _T_28639 & 10'h200;
  assign _T_28642 = _T_28640 == 10'h0;
  assign _T_28648 = _T_25900 ^ 10'h1c7;
  assign _T_28649 = _T_28648 & 10'h200;
  assign _T_28651 = _T_28649 == 10'h0;
  assign _T_28657 = _T_25900 ^ 10'hdf;
  assign _T_28658 = _T_28657 & 10'h200;
  assign _T_28660 = _T_28658 == 10'h0;
  assign _T_28666 = _T_25900 ^ 10'h18a;
  assign _T_28667 = _T_28666 & 10'h200;
  assign _T_28669 = _T_28667 == 10'h0;
  assign _T_28675 = _T_25900 ^ 10'h132;
  assign _T_28676 = _T_28675 & 10'h200;
  assign _T_28678 = _T_28676 == 10'h0;
  assign _T_28684 = _T_25900 ^ 10'h12b;
  assign _T_28685 = _T_28684 & 10'h200;
  assign _T_28687 = _T_28685 == 10'h0;
  assign _T_28693 = _T_25900 ^ 10'h10b;
  assign _T_28694 = _T_28693 & 10'h200;
  assign _T_28696 = _T_28694 == 10'h0;
  assign _T_28702 = _T_25900 ^ 10'h1f9;
  assign _T_28703 = _T_28702 & 10'h200;
  assign _T_28705 = _T_28703 == 10'h0;
  assign _T_28711 = _T_25900 ^ 10'h1b6;
  assign _T_28712 = _T_28711 & 10'h200;
  assign _T_28714 = _T_28712 == 10'h0;
  assign _T_28720 = _T_25900 ^ 10'h1af;
  assign _T_28721 = _T_28720 & 10'h200;
  assign _T_28723 = _T_28721 == 10'h0;
  assign _T_28729 = _T_25900 ^ 10'h1d9;
  assign _T_28730 = _T_28729 & 10'h200;
  assign _T_28732 = _T_28730 == 10'h0;
  assign _T_28738 = _T_25900 ^ 10'h1ea;
  assign _T_28739 = _T_28738 & 10'h200;
  assign _T_28741 = _T_28739 == 10'h0;
  assign _T_28747 = _T_25900 ^ 10'h1aa;
  assign _T_28748 = _T_28747 & 10'h200;
  assign _T_28750 = _T_28748 == 10'h0;
  assign _T_28756 = _T_25900 ^ 10'h213;
  assign _T_28757 = _T_28756 & 10'h200;
  assign _T_28759 = _T_28757 == 10'h0;
  assign _T_28765 = _T_25900 ^ 10'h176;
  assign _T_28766 = _T_28765 & 10'h200;
  assign _T_28768 = _T_28766 == 10'h0;
  assign _T_28774 = _T_25900 ^ 10'hd1;
  assign _T_28775 = _T_28774 & 10'h200;
  assign _T_28777 = _T_28775 == 10'h0;
  assign _T_28783 = _T_25900 ^ 10'h1e7;
  assign _T_28784 = _T_28783 & 10'h200;
  assign _T_28786 = _T_28784 == 10'h0;
  assign _T_28792 = _T_25900 ^ 10'h204;
  assign _T_28793 = _T_28792 & 10'h200;
  assign _T_28795 = _T_28793 == 10'h0;
  assign _T_28801 = _T_25900 ^ 10'h156;
  assign _T_28802 = _T_28801 & 10'h200;
  assign _T_28804 = _T_28802 == 10'h0;
  assign _T_28810 = _T_25900 ^ 10'h163;
  assign _T_28811 = _T_28810 & 10'h200;
  assign _T_28813 = _T_28811 == 10'h0;
  assign _T_28819 = _T_25900 ^ 10'h1ca;
  assign _T_28820 = _T_28819 & 10'h200;
  assign _T_28822 = _T_28820 == 10'h0;
  assign _T_28828 = _T_25900 ^ 10'h20d;
  assign _T_28829 = _T_28828 & 10'h200;
  assign _T_28831 = _T_28829 == 10'h0;
  assign _T_28837 = _T_25900 ^ 10'h127;
  assign _T_28838 = _T_28837 & 10'h200;
  assign _T_28840 = _T_28838 == 10'h0;
  assign _T_28846 = _T_25900 ^ 10'h11a;
  assign _T_28847 = _T_28846 & 10'h200;
  assign _T_28849 = _T_28847 == 10'h0;
  assign _T_28855 = _T_25900 ^ 10'h19e;
  assign _T_28856 = _T_28855 & 10'h200;
  assign _T_28858 = _T_28856 == 10'h0;
  assign _T_28864 = _T_25900 ^ 10'h147;
  assign _T_28865 = _T_28864 & 10'h200;
  assign _T_28867 = _T_28865 == 10'h0;
  assign _T_28873 = _T_25900 ^ 10'h199;
  assign _T_28874 = _T_28873 & 10'h200;
  assign _T_28876 = _T_28874 == 10'h0;
  assign _T_28882 = _T_25900 ^ 10'h107;
  assign _T_28883 = _T_28882 & 10'h200;
  assign _T_28885 = _T_28883 == 10'h0;
  assign _T_28891 = _T_25900 ^ 10'h136;
  assign _T_28892 = _T_28891 & 10'h200;
  assign _T_28894 = _T_28892 == 10'h0;
  assign _T_28900 = _T_25900 ^ 10'h43;
  assign _T_28901 = _T_28900 & 10'h200;
  assign _T_28903 = _T_28901 == 10'h0;
  assign _T_28909 = _T_25900 ^ 10'h14b;
  assign _T_28910 = _T_28909 & 10'h200;
  assign _T_28912 = _T_28910 == 10'h0;
  assign _T_28918 = _T_25900 ^ 10'h1b9;
  assign _T_28919 = _T_28918 & 10'h200;
  assign _T_28921 = _T_28919 == 10'h0;
  assign _T_28927 = _T_25900 ^ 10'h172;
  assign _T_28928 = _T_28927 & 10'h200;
  assign _T_28930 = _T_28928 == 10'h0;
  assign _T_28936 = _T_25900 ^ 10'h1f6;
  assign _T_28937 = _T_28936 & 10'h200;
  assign _T_28939 = _T_28937 == 10'h0;
  assign _T_28945 = _T_25900 ^ 10'h1cf;
  assign _T_28946 = _T_28945 & 10'h200;
  assign _T_28948 = _T_28946 == 10'h0;
  assign _T_28954 = _T_25900 ^ 10'h152;
  assign _T_28955 = _T_28954 & 10'h200;
  assign _T_28957 = _T_28955 == 10'h0;
  assign _T_28963 = _T_25900 ^ 10'h1d6;
  assign _T_28964 = _T_28963 & 10'h200;
  assign _T_28966 = _T_28964 == 10'h0;
  assign _T_28972 = _T_25900 ^ 10'h167;
  assign _T_28973 = _T_28972 & 10'h200;
  assign _T_28975 = _T_28973 == 10'h0;
  assign _T_28981 = _T_25900 ^ 10'h150;
  assign _T_28982 = _T_28981 & 10'h200;
  assign _T_28984 = _T_28982 == 10'h0;
  assign _T_28990 = _T_25900 ^ 10'h182;
  assign _T_28991 = _T_28990 & 10'h200;
  assign _T_28993 = _T_28991 == 10'h0;
  assign _T_28999 = _T_25900 ^ 10'h13a;
  assign _T_29000 = _T_28999 & 10'h200;
  assign _T_29002 = _T_29000 == 10'h0;
  assign _T_29008 = _T_25900 ^ 10'h1be;
  assign _T_29009 = _T_29008 & 10'h200;
  assign _T_29011 = _T_29009 == 10'h0;
  assign _T_29017 = _T_25900 ^ 10'h1f1;
  assign _T_29018 = _T_29017 & 10'h200;
  assign _T_29020 = _T_29018 == 10'h0;
  assign _T_29026 = _T_25900 ^ 10'h1d1;
  assign _T_29027 = _T_29026 & 10'h200;
  assign _T_29029 = _T_29027 == 10'h0;
  assign _T_29035 = _T_25900 ^ 10'h1c2;
  assign _T_29036 = _T_29035 & 10'h200;
  assign _T_29038 = _T_29036 == 10'h0;
  assign _T_29044 = _T_25900 ^ 10'h16b;
  assign _T_29045 = _T_29044 & 10'h200;
  assign _T_29047 = _T_29045 == 10'h0;
  assign _T_29053 = _T_25900 ^ 10'h1e2;
  assign _T_29054 = _T_29053 & 10'h200;
  assign _T_29056 = _T_29054 == 10'h0;
  assign _T_29062 = _T_25900 ^ 10'h20c;
  assign _T_29063 = _T_29062 & 10'h200;
  assign _T_29065 = _T_29063 == 10'h0;
  assign _T_29071 = _T_25900 ^ 10'h1ef;
  assign _T_29072 = _T_29071 & 10'h200;
  assign _T_29074 = _T_29072 == 10'h0;
  assign _T_29080 = _T_25900 ^ 10'hda;
  assign _T_29081 = _T_29080 & 10'h200;
  assign _T_29083 = _T_29081 == 10'h0;
  assign _T_29089 = _T_25900 ^ 10'h170;
  assign _T_29090 = _T_29089 & 10'h200;
  assign _T_29092 = _T_29090 == 10'h0;
  assign _T_29098 = _T_25900 ^ 10'h205;
  assign _T_29099 = _T_29098 & 10'h200;
  assign _T_29101 = _T_29099 == 10'h0;
  assign _T_29107 = _T_25900 ^ 10'h13f;
  assign _T_29108 = _T_29107 & 10'h200;
  assign _T_29110 = _T_29108 == 10'h0;
  assign _T_29116 = _T_25900 ^ 10'h130;
  assign _T_29117 = _T_29116 & 10'h200;
  assign _T_29119 = _T_29117 == 10'h0;
  assign _T_29125 = _T_25900 ^ 10'h102;
  assign _T_29126 = _T_29125 & 10'h200;
  assign _T_29128 = _T_29126 == 10'h0;
  assign _T_29134 = _T_25900 ^ 10'h15f;
  assign _T_29135 = _T_29134 & 10'h200;
  assign _T_29137 = _T_29135 == 10'h0;
  assign _T_29143 = _T_25900 ^ 10'h186;
  assign _T_29144 = _T_29143 & 10'h200;
  assign _T_29146 = _T_29144 == 10'h0;
  assign _T_29152 = _T_25900 ^ 10'h191;
  assign _T_29153 = _T_29152 & 10'h200;
  assign _T_29155 = _T_29153 == 10'h0;
  assign _T_29161 = _T_25900 ^ 10'h1a2;
  assign _T_29162 = _T_29161 & 10'h200;
  assign _T_29164 = _T_29162 == 10'h0;
  assign _T_29170 = _T_25900 ^ 10'h122;
  assign _T_29171 = _T_29170 & 10'h200;
  assign _T_29173 = _T_29171 == 10'h0;
  assign _T_29179 = _T_25900 ^ 10'h17a;
  assign _T_29180 = _T_29179 & 10'h200;
  assign _T_29182 = _T_29180 == 10'h0;
  assign _T_29188 = _T_25900 ^ 10'h1b1;
  assign _T_29189 = _T_29188 & 10'h200;
  assign _T_29191 = _T_29189 == 10'h0;
  assign _T_29197 = _T_25900 ^ 10'h1fe;
  assign _T_29198 = _T_29197 & 10'h200;
  assign _T_29200 = _T_29198 == 10'h0;
  assign _T_29206 = _T_25900 ^ 10'hcf;
  assign _T_29207 = _T_29206 & 10'h200;
  assign _T_29209 = _T_29207 == 10'h0;
  assign _T_29215 = _T_25900 ^ 10'h1de;
  assign _T_29216 = _T_29215 & 10'h200;
  assign _T_29218 = _T_29216 == 10'h0;
  assign _T_29224 = _T_25900 ^ 10'h110;
  assign _T_29225 = _T_29224 & 10'h200;
  assign _T_29227 = _T_29225 == 10'h0;
  assign _T_29233 = _T_25900 ^ 10'h17f;
  assign _T_29234 = _T_29233 & 10'h200;
  assign _T_29236 = _T_29234 == 10'h0;
  assign _T_29242 = _T_25900 ^ 10'h15a;
  assign _T_29243 = _T_29242 & 10'h200;
  assign _T_29245 = _T_29243 == 10'h0;
  assign _T_29251 = _T_25900 ^ 10'hd6;
  assign _T_29252 = _T_29251 & 10'h200;
  assign _T_29254 = _T_29252 == 10'h0;
  assign _T_29260 = _T_25900 ^ 10'h11f;
  assign _T_29261 = _T_29260 & 10'h200;
  assign _T_29263 = _T_29261 == 10'h0;
  assign _T_29269 = _T_25900 ^ 10'h12c;
  assign _T_29270 = _T_29269 & 10'h200;
  assign _T_29272 = _T_29270 == 10'h0;
  assign _T_29278 = _T_25900 ^ 10'h1bf;
  assign _T_29279 = _T_29278 & 10'h200;
  assign _T_29281 = _T_29279 == 10'h0;
  assign _T_29287 = _T_25900 ^ 10'h13b;
  assign _T_29288 = _T_29287 & 10'h200;
  assign _T_29290 = _T_29288 == 10'h0;
  assign _T_29296 = _T_25900 ^ 10'h1b0;
  assign _T_29297 = _T_29296 & 10'h200;
  assign _T_29299 = _T_29297 == 10'h0;
  assign _T_29305 = _T_25900 ^ 10'h19a;
  assign _T_29306 = _T_29305 & 10'h200;
  assign _T_29308 = _T_29306 == 10'h0;
  assign _T_29314 = _T_25900 ^ 10'h106;
  assign _T_29315 = _T_29314 & 10'h200;
  assign _T_29317 = _T_29315 == 10'h0;
  assign _T_29323 = _T_25900 ^ 10'h195;
  assign _T_29324 = _T_29323 & 10'h200;
  assign _T_29326 = _T_29324 == 10'h0;
  assign _T_29332 = _T_25900 ^ 10'h1a6;
  assign _T_29333 = _T_29332 & 10'h200;
  assign _T_29335 = _T_29333 == 10'h0;
  assign _T_29341 = _T_25900 ^ 10'h111;
  assign _T_29342 = _T_29341 & 10'h200;
  assign _T_29344 = _T_29342 == 10'h0;
  assign _T_29350 = _T_25900 ^ 10'h175;
  assign _T_29351 = _T_29350 & 10'h200;
  assign _T_29353 = _T_29351 == 10'h0;
  assign _T_29359 = _T_25900 ^ 10'h131;
  assign _T_29360 = _T_29359 & 10'h200;
  assign _T_29362 = _T_29360 == 10'h0;
  assign _T_29368 = _T_25900 ^ 10'hd2;
  assign _T_29369 = _T_29368 & 10'h200;
  assign _T_29371 = _T_29369 == 10'h0;
  assign _T_29377 = _T_25900 ^ 10'h146;
  assign _T_29378 = _T_29377 & 10'h200;
  assign _T_29380 = _T_29378 == 10'h0;
  assign _T_29386 = _T_25900 ^ 10'h126;
  assign _T_29387 = _T_29386 & 10'h200;
  assign _T_29389 = _T_29387 == 10'h0;
  assign _T_29395 = _T_25900 ^ 10'h155;
  assign _T_29396 = _T_29395 & 10'h200;
  assign _T_29398 = _T_29396 == 10'h0;
  assign _T_29404 = _T_25900 ^ 10'h1fa;
  assign _T_29405 = _T_29404 & 10'h200;
  assign _T_29407 = _T_29405 == 10'h0;
  assign _T_29413 = _T_25900 ^ 10'h10c;
  assign _T_29414 = _T_29413 & 10'h200;
  assign _T_29416 = _T_29414 == 10'h0;
  assign _T_29422 = _T_25900 ^ 10'h166;
  assign _T_29423 = _T_29422 & 10'h200;
  assign _T_29425 = _T_29423 == 10'h0;
  assign _T_29431 = _T_25900 ^ 10'h1b5;
  assign _T_29432 = _T_29431 & 10'h200;
  assign _T_29434 = _T_29432 == 10'h0;
  assign _T_29440 = _T_25900 ^ 10'h1da;
  assign _T_29441 = _T_29440 & 10'h200;
  assign _T_29443 = _T_29441 == 10'h0;
  assign _T_29449 = _T_25900 ^ 10'h190;
  assign _T_29450 = _T_29449 & 10'h200;
  assign _T_29452 = _T_29450 == 10'h0;
  assign _T_29458 = _T_25900 ^ 10'h214;
  assign _T_29459 = _T_29458 & 10'h200;
  assign _T_29461 = _T_29459 == 10'h0;
  assign _T_29467 = _T_25900 ^ 10'h11b;
  assign _T_29468 = _T_29467 & 10'h200;
  assign _T_29470 = _T_29468 == 10'h0;
  assign _T_29476 = _T_25900 ^ 10'h19f;
  assign _T_29477 = _T_29476 & 10'h200;
  assign _T_29479 = _T_29477 == 10'h0;
  assign _T_29485 = _T_25900 ^ 10'h18b;
  assign _T_29486 = _T_29485 & 10'h200;
  assign _T_29488 = _T_29486 == 10'h0;
  assign _T_29494 = _T_25900 ^ 10'h1d0;
  assign _T_29495 = _T_29494 & 10'h200;
  assign _T_29497 = _T_29495 == 10'h0;
  assign _T_29503 = _T_25900 ^ 10'h14c;
  assign _T_29504 = _T_29503 & 10'h200;
  assign _T_29506 = _T_29504 == 10'h0;
  assign _T_29512 = _T_25900 ^ 10'h1ab;
  assign _T_29513 = _T_29512 & 10'h200;
  assign _T_29515 = _T_29513 == 10'h0;
  assign _T_29521 = _T_25900 ^ 10'h210;
  assign _T_29522 = _T_29521 & 10'h200;
  assign _T_29524 = _T_29522 == 10'h0;
  assign _T_29530 = _T_25900 ^ 10'h1cb;
  assign _T_29531 = _T_29530 & 10'h200;
  assign _T_29533 = _T_29531 == 10'h0;
  assign _T_29539 = _T_25900 ^ 10'h115;
  assign _T_29540 = _T_29539 & 10'h200;
  assign _T_29542 = _T_29540 == 10'h0;
  assign _T_29548 = _T_25900 ^ 10'h1ba;
  assign _T_29549 = _T_29548 & 10'h200;
  assign _T_29551 = _T_29549 == 10'h0;
  assign _T_29557 = _T_25900 ^ 10'h1f5;
  assign _T_29558 = _T_29557 & 10'h200;
  assign _T_29560 = _T_29558 == 10'h0;
  assign _T_29566 = _T_25900 ^ 10'h171;
  assign _T_29567 = _T_29566 & 10'h200;
  assign _T_29569 = _T_29567 == 10'h0;
  assign _T_29575 = _T_25900 ^ 10'h142;
  assign _T_29576 = _T_29575 & 10'h200;
  assign _T_29578 = _T_29576 == 10'h0;
  assign _T_29584 = _T_25900 ^ 10'h1e6;
  assign _T_29585 = _T_29584 & 10'h200;
  assign _T_29587 = _T_29585 == 10'h0;
  assign _T_29593 = _T_25900 ^ 10'h151;
  assign _T_29594 = _T_29593 & 10'h200;
  assign _T_29596 = _T_29594 == 10'h0;
  assign _T_29602 = _T_25900 ^ 10'h1d5;
  assign _T_29603 = _T_29602 & 10'h200;
  assign _T_29605 = _T_29603 == 10'h0;
  assign _T_29611 = _T_25900 ^ 10'h162;
  assign _T_29612 = _T_29611 & 10'h200;
  assign _T_29614 = _T_29612 == 10'h0;
  assign _T_29620 = _T_25900 ^ 10'h135;
  assign _T_29621 = _T_29620 & 10'h200;
  assign _T_29623 = _T_29621 == 10'h0;
  assign _T_29629 = _T_25900 ^ 10'hd7;
  assign _T_29630 = _T_29629 & 10'h200;
  assign _T_29632 = _T_29630 == 10'h0;
  assign _T_29638 = _T_25900 ^ 10'h1eb;
  assign _T_29639 = _T_29638 & 10'h200;
  assign _T_29641 = _T_29639 == 10'h0;
  assign _T_29647 = _T_25900 ^ 10'hde;
  assign _T_29648 = _T_29647 & 10'h200;
  assign _T_29650 = _T_29648 == 10'h0;
  assign _T_29656 = _T_25900 ^ 10'h1f0;
  assign _T_29657 = _T_29656 & 10'h200;
  assign _T_29659 = _T_29657 == 10'h0;
  assign _T_29665 = _T_25900 ^ 10'h1c6;
  assign _T_29666 = _T_29665 & 10'h200;
  assign _T_29668 = _T_29666 == 10'h0;
  assign _T_29674 = _T_25900 ^ 10'h16c;
  assign _T_29675 = _T_29674 & 10'h200;
  assign _T_29677 = _T_29675 == 10'h0;
  assign _T_34998 = io_hart_in_0_a_bits_mask[0];
  assign _T_34999 = io_hart_in_0_a_bits_mask[1];
  assign _T_35000 = io_hart_in_0_a_bits_mask[2];
  assign _T_35001 = io_hart_in_0_a_bits_mask[3];
  assign _T_35005 = _T_34998 ? 8'hff : 8'h0;
  assign _T_35009 = _T_34999 ? 8'hff : 8'h0;
  assign _T_35013 = _T_35000 ? 8'hff : 8'h0;
  assign _T_35017 = _T_35001 ? 8'hff : 8'h0;
  assign _T_35018 = {_T_35009,_T_35005};
  assign _T_35019 = {_T_35017,_T_35013};
  assign _T_35020 = {_T_35019,_T_35018};
  assign _T_35044 = _T_35020[7:0];
  assign _T_35048 = ~ _T_35044;
  assign _T_35050 = _T_35048 == 8'h0;
  assign _T_35064 = io_hart_in_0_a_bits_data[7:0];
  assign _T_35084 = _T_35020[15:8];
  assign _T_35088 = ~ _T_35084;
  assign _T_35090 = _T_35088 == 8'h0;
  assign _T_35104 = io_hart_in_0_a_bits_data[15:8];
  assign _GEN_5773 = {{8'd0}, _T_24620};
  assign _T_35119 = _GEN_5773 << 8;
  assign _GEN_5774 = {{8'd0}, _T_24618};
  assign _T_35123 = _GEN_5774 | _T_35119;
  assign _T_35124 = _T_35020[23:16];
  assign _T_35128 = ~ _T_35124;
  assign _T_35130 = _T_35128 == 8'h0;
  assign _T_35144 = io_hart_in_0_a_bits_data[23:16];
  assign _GEN_5775 = {{16'd0}, _T_24622};
  assign _T_35159 = _GEN_5775 << 16;
  assign _GEN_5776 = {{8'd0}, _T_35123};
  assign _T_35163 = _GEN_5776 | _T_35159;
  assign _T_35164 = _T_35020[31:24];
  assign _T_35168 = ~ _T_35164;
  assign _T_35170 = _T_35168 == 8'h0;
  assign _T_35184 = io_hart_in_0_a_bits_data[31:24];
  assign _GEN_5777 = {{24'd0}, _T_24624};
  assign _T_35199 = _GEN_5777 << 24;
  assign _GEN_5778 = {{8'd0}, _T_35163};
  assign _T_35203 = _GEN_5778 | _T_35199;
  assign _GEN_5779 = {{8'd0}, _T_25532};
  assign _T_35279 = _GEN_5779 << 8;
  assign _GEN_5780 = {{8'd0}, _T_25530};
  assign _T_35283 = _GEN_5780 | _T_35279;
  assign _GEN_5781 = {{16'd0}, _T_25534};
  assign _T_35319 = _GEN_5781 << 16;
  assign _GEN_5782 = {{8'd0}, _T_35283};
  assign _T_35323 = _GEN_5782 | _T_35319;
  assign _GEN_5783 = {{24'd0}, _T_25536};
  assign _T_35359 = _GEN_5783 << 24;
  assign _GEN_5784 = {{8'd0}, _T_35323};
  assign _T_35363 = _GEN_5784 | _T_35359;
  assign _GEN_5785 = {{8'd0}, _T_24476};
  assign _T_35439 = _GEN_5785 << 8;
  assign _GEN_5786 = {{8'd0}, _T_24474};
  assign _T_35443 = _GEN_5786 | _T_35439;
  assign _GEN_5787 = {{16'd0}, _T_24478};
  assign _T_35479 = _GEN_5787 << 16;
  assign _GEN_5788 = {{8'd0}, _T_35443};
  assign _T_35483 = _GEN_5788 | _T_35479;
  assign _GEN_5789 = {{24'd0}, _T_24480};
  assign _T_35519 = _GEN_5789 << 24;
  assign _GEN_5790 = {{8'd0}, _T_35483};
  assign _T_35523 = _GEN_5790 | _T_35519;
  assign _GEN_5791 = {{8'd0}, _T_24364};
  assign _T_35599 = _GEN_5791 << 8;
  assign _GEN_5792 = {{8'd0}, _T_24362};
  assign _T_35603 = _GEN_5792 | _T_35599;
  assign _GEN_5793 = {{16'd0}, _T_24366};
  assign _T_35639 = _GEN_5793 << 16;
  assign _GEN_5794 = {{8'd0}, _T_35603};
  assign _T_35643 = _GEN_5794 | _T_35639;
  assign _GEN_5795 = {{24'd0}, _T_24368};
  assign _T_35679 = _GEN_5795 << 24;
  assign _GEN_5796 = {{8'd0}, _T_35643};
  assign _T_35683 = _GEN_5796 | _T_35679;
  assign _GEN_5797 = {{8'd0}, _T_25444};
  assign _T_35919 = _GEN_5797 << 8;
  assign _GEN_5798 = {{8'd0}, _T_25442};
  assign _T_35923 = _GEN_5798 | _T_35919;
  assign _GEN_5799 = {{16'd0}, _T_25446};
  assign _T_35959 = _GEN_5799 << 16;
  assign _GEN_5800 = {{8'd0}, _T_35923};
  assign _T_35963 = _GEN_5800 | _T_35959;
  assign _GEN_5801 = {{24'd0}, _T_25448};
  assign _T_35999 = _GEN_5801 << 24;
  assign _GEN_5802 = {{8'd0}, _T_35963};
  assign _T_36003 = _GEN_5802 | _T_35999;
  assign _GEN_5803 = {{8'd0}, _T_25548};
  assign _T_36079 = _GEN_5803 << 8;
  assign _GEN_5804 = {{8'd0}, _T_25546};
  assign _T_36083 = _GEN_5804 | _T_36079;
  assign _GEN_5805 = {{16'd0}, _T_25550};
  assign _T_36119 = _GEN_5805 << 16;
  assign _GEN_5806 = {{8'd0}, _T_36083};
  assign _T_36123 = _GEN_5806 | _T_36119;
  assign _GEN_5807 = {{24'd0}, _T_25552};
  assign _T_36159 = _GEN_5807 << 24;
  assign _GEN_5808 = {{8'd0}, _T_36123};
  assign _T_36163 = _GEN_5808 | _T_36159;
  assign _GEN_5809 = {{8'd0}, _T_24516};
  assign _T_36239 = _GEN_5809 << 8;
  assign _GEN_5810 = {{8'd0}, _T_24514};
  assign _T_36243 = _GEN_5810 | _T_36239;
  assign _GEN_5811 = {{16'd0}, _T_24518};
  assign _T_36279 = _GEN_5811 << 16;
  assign _GEN_5812 = {{8'd0}, _T_36243};
  assign _T_36283 = _GEN_5812 | _T_36279;
  assign _GEN_5813 = {{24'd0}, _T_24520};
  assign _T_36319 = _GEN_5813 << 24;
  assign _GEN_5814 = {{8'd0}, _T_36283};
  assign _T_36323 = _GEN_5814 | _T_36319;
  assign _GEN_5815 = {{8'd0}, _T_24964};
  assign _T_36399 = _GEN_5815 << 8;
  assign _GEN_5816 = {{8'd0}, _T_24962};
  assign _T_36403 = _GEN_5816 | _T_36399;
  assign _GEN_5817 = {{16'd0}, _T_24966};
  assign _T_36439 = _GEN_5817 << 16;
  assign _GEN_5818 = {{8'd0}, _T_36403};
  assign _T_36443 = _GEN_5818 | _T_36439;
  assign _GEN_5819 = {{24'd0}, _T_24968};
  assign _T_36479 = _GEN_5819 << 24;
  assign _GEN_5820 = {{8'd0}, _T_36443};
  assign _T_36483 = _GEN_5820 | _T_36479;
  assign _T_36663 = _T_99498 & _T_35050;
  assign _GEN_2439 = _T_36663 ? _T_35064 : _GEN_357;
  assign _T_36703 = _T_99498 & _T_35090;
  assign _GEN_2440 = _T_36703 ? _T_35104 : _GEN_358;
  assign _T_36743 = _T_99498 & _T_35130;
  assign _GEN_2441 = _T_36743 ? _T_35144 : _GEN_359;
  assign _T_36783 = _T_99498 & _T_35170;
  assign _GEN_2442 = _T_36783 ? _T_35184 : _GEN_360;
  assign _GEN_5827 = {{8'd0}, _T_23908};
  assign _T_36879 = _GEN_5827 << 8;
  assign _GEN_5828 = {{8'd0}, _T_23906};
  assign _T_36883 = _GEN_5828 | _T_36879;
  assign _GEN_5829 = {{16'd0}, _T_23910};
  assign _T_36919 = _GEN_5829 << 16;
  assign _GEN_5830 = {{8'd0}, _T_36883};
  assign _T_36923 = _GEN_5830 | _T_36919;
  assign _GEN_5831 = {{24'd0}, _T_23912};
  assign _T_36959 = _GEN_5831 << 24;
  assign _GEN_5832 = {{8'd0}, _T_36923};
  assign _T_36963 = _GEN_5832 | _T_36959;
  assign _GEN_5833 = {{8'd0}, _T_24164};
  assign _T_37039 = _GEN_5833 << 8;
  assign _GEN_5834 = {{8'd0}, _T_24162};
  assign _T_37043 = _GEN_5834 | _T_37039;
  assign _GEN_5835 = {{16'd0}, _T_24166};
  assign _T_37079 = _GEN_5835 << 16;
  assign _GEN_5836 = {{8'd0}, _T_37043};
  assign _T_37083 = _GEN_5836 | _T_37079;
  assign _GEN_5837 = {{24'd0}, _T_24168};
  assign _T_37119 = _GEN_5837 << 24;
  assign _GEN_5838 = {{8'd0}, _T_37083};
  assign _T_37123 = _GEN_5838 | _T_37119;
  assign _GEN_5839 = {{8'd0}, _T_25292};
  assign _T_37199 = _GEN_5839 << 8;
  assign _GEN_5840 = {{8'd0}, _T_25290};
  assign _T_37203 = _GEN_5840 | _T_37199;
  assign _GEN_5841 = {{16'd0}, _T_25294};
  assign _T_37239 = _GEN_5841 << 16;
  assign _GEN_5842 = {{8'd0}, _T_37203};
  assign _T_37243 = _GEN_5842 | _T_37239;
  assign _GEN_5843 = {{24'd0}, _T_25296};
  assign _T_37279 = _GEN_5843 << 24;
  assign _GEN_5844 = {{8'd0}, _T_37243};
  assign _T_37283 = _GEN_5844 | _T_37279;
  assign _GEN_5845 = {{8'd0}, _T_24732};
  assign _T_37359 = _GEN_5845 << 8;
  assign _GEN_5846 = {{8'd0}, _T_24730};
  assign _T_37363 = _GEN_5846 | _T_37359;
  assign _GEN_5847 = {{16'd0}, _T_24734};
  assign _T_37399 = _GEN_5847 << 16;
  assign _GEN_5848 = {{8'd0}, _T_37363};
  assign _T_37403 = _GEN_5848 | _T_37399;
  assign _GEN_5849 = {{24'd0}, _T_24736};
  assign _T_37439 = _GEN_5849 << 24;
  assign _GEN_5850 = {{8'd0}, _T_37403};
  assign _T_37443 = _GEN_5850 | _T_37439;
  assign _GEN_5851 = {{8'd0}, _T_25220};
  assign _T_37519 = _GEN_5851 << 8;
  assign _GEN_5852 = {{8'd0}, _T_25218};
  assign _T_37523 = _GEN_5852 | _T_37519;
  assign _GEN_5853 = {{16'd0}, _T_25222};
  assign _T_37559 = _GEN_5853 << 16;
  assign _GEN_5854 = {{8'd0}, _T_37523};
  assign _T_37563 = _GEN_5854 | _T_37559;
  assign _GEN_5855 = {{24'd0}, _T_25224};
  assign _T_37599 = _GEN_5855 << 24;
  assign _GEN_5856 = {{8'd0}, _T_37563};
  assign _T_37603 = _GEN_5856 | _T_37599;
  assign _GEN_5857 = {{8'd0}, _T_25788};
  assign _T_37679 = _GEN_5857 << 8;
  assign _GEN_5858 = {{8'd0}, _T_25786};
  assign _T_37683 = _GEN_5858 | _T_37679;
  assign _GEN_5859 = {{16'd0}, _T_25790};
  assign _T_37719 = _GEN_5859 << 16;
  assign _GEN_5860 = {{8'd0}, _T_37683};
  assign _T_37723 = _GEN_5860 | _T_37719;
  assign _GEN_5861 = {{24'd0}, _T_25792};
  assign _T_37759 = _GEN_5861 << 24;
  assign _GEN_5862 = {{8'd0}, _T_37723};
  assign _T_37763 = _GEN_5862 | _T_37759;
  assign _GEN_5863 = {{8'd0}, _T_23852};
  assign _T_37839 = _GEN_5863 << 8;
  assign _GEN_5864 = {{8'd0}, _T_23850};
  assign _T_37843 = _GEN_5864 | _T_37839;
  assign _GEN_5865 = {{16'd0}, _T_23854};
  assign _T_37879 = _GEN_5865 << 16;
  assign _GEN_5866 = {{8'd0}, _T_37843};
  assign _T_37883 = _GEN_5866 | _T_37879;
  assign _GEN_5867 = {{24'd0}, _T_23856};
  assign _T_37919 = _GEN_5867 << 24;
  assign _GEN_5868 = {{8'd0}, _T_37883};
  assign _T_37923 = _GEN_5868 | _T_37919;
  assign _GEN_5869 = {{8'd0}, _T_24780};
  assign _T_37999 = _GEN_5869 << 8;
  assign _GEN_5870 = {{8'd0}, _T_24778};
  assign _T_38003 = _GEN_5870 | _T_37999;
  assign _GEN_5871 = {{16'd0}, _T_24782};
  assign _T_38039 = _GEN_5871 << 16;
  assign _GEN_5872 = {{8'd0}, _T_38003};
  assign _T_38043 = _GEN_5872 | _T_38039;
  assign _GEN_5873 = {{24'd0}, _T_24784};
  assign _T_38079 = _GEN_5873 << 24;
  assign _GEN_5874 = {{8'd0}, _T_38043};
  assign _T_38083 = _GEN_5874 | _T_38079;
  assign _GEN_5875 = {{8'd0}, _T_24772};
  assign _T_38159 = _GEN_5875 << 8;
  assign _GEN_5876 = {{8'd0}, _T_24770};
  assign _T_38163 = _GEN_5876 | _T_38159;
  assign _GEN_5877 = {{16'd0}, _T_24774};
  assign _T_38199 = _GEN_5877 << 16;
  assign _GEN_5878 = {{8'd0}, _T_38163};
  assign _T_38203 = _GEN_5878 | _T_38199;
  assign _GEN_5879 = {{24'd0}, _T_24776};
  assign _T_38239 = _GEN_5879 << 24;
  assign _GEN_5880 = {{8'd0}, _T_38203};
  assign _T_38243 = _GEN_5880 | _T_38239;
  assign _GEN_5881 = {{8'd0}, _T_25700};
  assign _T_38479 = _GEN_5881 << 8;
  assign _GEN_5882 = {{8'd0}, _T_25698};
  assign _T_38483 = _GEN_5882 | _T_38479;
  assign _GEN_5883 = {{16'd0}, _T_25702};
  assign _T_38519 = _GEN_5883 << 16;
  assign _GEN_5884 = {{8'd0}, _T_38483};
  assign _T_38523 = _GEN_5884 | _T_38519;
  assign _GEN_5885 = {{24'd0}, _T_25704};
  assign _T_38559 = _GEN_5885 << 24;
  assign _GEN_5886 = {{8'd0}, _T_38523};
  assign _T_38563 = _GEN_5886 | _T_38559;
  assign _GEN_5887 = {{8'd0}, _T_25476};
  assign _T_38639 = _GEN_5887 << 8;
  assign _GEN_5888 = {{8'd0}, _T_25474};
  assign _T_38643 = _GEN_5888 | _T_38639;
  assign _GEN_5889 = {{16'd0}, _T_25478};
  assign _T_38679 = _GEN_5889 << 16;
  assign _GEN_5890 = {{8'd0}, _T_38643};
  assign _T_38683 = _GEN_5890 | _T_38679;
  assign _GEN_5891 = {{24'd0}, _T_25480};
  assign _T_38719 = _GEN_5891 << 24;
  assign _GEN_5892 = {{8'd0}, _T_38683};
  assign _T_38723 = _GEN_5892 | _T_38719;
  assign _GEN_5893 = {{8'd0}, _T_24420};
  assign _T_38799 = _GEN_5893 << 8;
  assign _GEN_5894 = {{8'd0}, _T_24418};
  assign _T_38803 = _GEN_5894 | _T_38799;
  assign _GEN_5895 = {{16'd0}, _T_24422};
  assign _T_38839 = _GEN_5895 << 16;
  assign _GEN_5896 = {{8'd0}, _T_38803};
  assign _T_38843 = _GEN_5896 | _T_38839;
  assign _GEN_5897 = {{24'd0}, _T_24424};
  assign _T_38879 = _GEN_5897 << 24;
  assign _GEN_5898 = {{8'd0}, _T_38843};
  assign _T_38883 = _GEN_5898 | _T_38879;
  assign _GEN_5899 = {{8'd0}, _T_24932};
  assign _T_38959 = _GEN_5899 << 8;
  assign _GEN_5900 = {{8'd0}, _T_24930};
  assign _T_38963 = _GEN_5900 | _T_38959;
  assign _GEN_5901 = {{16'd0}, _T_24934};
  assign _T_38999 = _GEN_5901 << 16;
  assign _GEN_5902 = {{8'd0}, _T_38963};
  assign _T_39003 = _GEN_5902 | _T_38999;
  assign _GEN_5903 = {{24'd0}, _T_24936};
  assign _T_39039 = _GEN_5903 << 24;
  assign _GEN_5904 = {{8'd0}, _T_39003};
  assign _T_39043 = _GEN_5904 | _T_39039;
  assign _GEN_5905 = {{8'd0}, _T_25036};
  assign _T_39119 = _GEN_5905 << 8;
  assign _GEN_5906 = {{8'd0}, _T_25034};
  assign _T_39123 = _GEN_5906 | _T_39119;
  assign _GEN_5907 = {{16'd0}, _T_25038};
  assign _T_39159 = _GEN_5907 << 16;
  assign _GEN_5908 = {{8'd0}, _T_39123};
  assign _T_39163 = _GEN_5908 | _T_39159;
  assign _GEN_5909 = {{24'd0}, _T_25040};
  assign _T_39199 = _GEN_5909 << 24;
  assign _GEN_5910 = {{8'd0}, _T_39163};
  assign _T_39203 = _GEN_5910 | _T_39199;
  assign _GEN_5911 = {{8'd0}, _T_24004};
  assign _T_39279 = _GEN_5911 << 8;
  assign _GEN_5912 = {{8'd0}, _T_24002};
  assign _T_39283 = _GEN_5912 | _T_39279;
  assign _GEN_5913 = {{16'd0}, _T_24006};
  assign _T_39319 = _GEN_5913 << 16;
  assign _GEN_5914 = {{8'd0}, _T_39283};
  assign _T_39323 = _GEN_5914 | _T_39319;
  assign _GEN_5915 = {{24'd0}, _T_24008};
  assign _T_39359 = _GEN_5915 << 24;
  assign _GEN_5916 = {{8'd0}, _T_39323};
  assign _T_39363 = _GEN_5916 | _T_39359;
  assign _GEN_5917 = {{8'd0}, _T_24108};
  assign _T_39439 = _GEN_5917 << 8;
  assign _GEN_5918 = {{8'd0}, _T_24106};
  assign _T_39443 = _GEN_5918 | _T_39439;
  assign _GEN_5919 = {{16'd0}, _T_24110};
  assign _T_39479 = _GEN_5919 << 16;
  assign _GEN_5920 = {{8'd0}, _T_39443};
  assign _T_39483 = _GEN_5920 | _T_39479;
  assign _GEN_5921 = {{24'd0}, _T_24112};
  assign _T_39519 = _GEN_5921 << 24;
  assign _GEN_5922 = {{8'd0}, _T_39483};
  assign _T_39523 = _GEN_5922 | _T_39519;
  assign _GEN_5923 = {{8'd0}, _T_24260};
  assign _T_39599 = _GEN_5923 << 8;
  assign _GEN_5924 = {{8'd0}, _T_24258};
  assign _T_39603 = _GEN_5924 | _T_39599;
  assign _GEN_5925 = {{16'd0}, _T_24262};
  assign _T_39639 = _GEN_5925 << 16;
  assign _GEN_5926 = {{8'd0}, _T_39603};
  assign _T_39643 = _GEN_5926 | _T_39639;
  assign _GEN_5927 = {{24'd0}, _T_24264};
  assign _T_39679 = _GEN_5927 << 24;
  assign _GEN_5928 = {{8'd0}, _T_39643};
  assign _T_39683 = _GEN_5928 | _T_39679;
  assign _GEN_5929 = {{8'd0}, _T_25188};
  assign _T_39759 = _GEN_5929 << 8;
  assign _GEN_5930 = {{8'd0}, _T_25186};
  assign _T_39763 = _GEN_5930 | _T_39759;
  assign _GEN_5931 = {{16'd0}, _T_25190};
  assign _T_39799 = _GEN_5931 << 16;
  assign _GEN_5932 = {{8'd0}, _T_39763};
  assign _T_39803 = _GEN_5932 | _T_39799;
  assign _GEN_5933 = {{24'd0}, _T_25192};
  assign _T_39839 = _GEN_5933 << 24;
  assign _GEN_5934 = {{8'd0}, _T_39803};
  assign _T_39843 = _GEN_5934 | _T_39839;
  assign _GEN_5935 = {{8'd0}, _T_23756};
  assign _T_39919 = _GEN_5935 << 8;
  assign _GEN_5936 = {{8'd0}, _T_23754};
  assign _T_39923 = _GEN_5936 | _T_39919;
  assign _GEN_5937 = {{16'd0}, _T_23758};
  assign _T_39959 = _GEN_5937 << 16;
  assign _GEN_5938 = {{8'd0}, _T_39923};
  assign _T_39963 = _GEN_5938 | _T_39959;
  assign _GEN_5939 = {{24'd0}, _T_23760};
  assign _T_39999 = _GEN_5939 << 24;
  assign _GEN_5940 = {{8'd0}, _T_39963};
  assign _T_40003 = _GEN_5940 | _T_39999;
  assign _GEN_5941 = {{8'd0}, _T_24812};
  assign _T_40079 = _GEN_5941 << 8;
  assign _GEN_5942 = {{8'd0}, _T_24810};
  assign _T_40083 = _GEN_5942 | _T_40079;
  assign _GEN_5943 = {{16'd0}, _T_24814};
  assign _T_40119 = _GEN_5943 << 16;
  assign _GEN_5944 = {{8'd0}, _T_40083};
  assign _T_40123 = _GEN_5944 | _T_40119;
  assign _GEN_5945 = {{24'd0}, _T_24816};
  assign _T_40159 = _GEN_5945 << 24;
  assign _GEN_5946 = {{8'd0}, _T_40123};
  assign _T_40163 = _GEN_5946 | _T_40159;
  assign _GEN_5947 = {{8'd0}, _T_24676};
  assign _T_40239 = _GEN_5947 << 8;
  assign _GEN_5948 = {{8'd0}, _T_24674};
  assign _T_40243 = _GEN_5948 | _T_40239;
  assign _GEN_5949 = {{16'd0}, _T_24678};
  assign _T_40279 = _GEN_5949 << 16;
  assign _GEN_5950 = {{8'd0}, _T_40243};
  assign _T_40283 = _GEN_5950 | _T_40279;
  assign _GEN_5951 = {{24'd0}, _T_24680};
  assign _T_40319 = _GEN_5951 << 24;
  assign _GEN_5952 = {{8'd0}, _T_40283};
  assign _T_40323 = _GEN_5952 | _T_40319;
  assign _GEN_5953 = {{8'd0}, _T_25732};
  assign _T_40399 = _GEN_5953 << 8;
  assign _GEN_5954 = {{8'd0}, _T_25730};
  assign _T_40403 = _GEN_5954 | _T_40399;
  assign _GEN_5955 = {{16'd0}, _T_25734};
  assign _T_40439 = _GEN_5955 << 16;
  assign _GEN_5956 = {{8'd0}, _T_40403};
  assign _T_40443 = _GEN_5956 | _T_40439;
  assign _GEN_5957 = {{24'd0}, _T_25736};
  assign _T_40479 = _GEN_5957 << 24;
  assign _GEN_5958 = {{8'd0}, _T_40443};
  assign _T_40483 = _GEN_5958 | _T_40479;
  assign _GEN_5959 = {{8'd0}, _T_24452};
  assign _T_40559 = _GEN_5959 << 8;
  assign _GEN_5960 = {{8'd0}, _T_24450};
  assign _T_40563 = _GEN_5960 | _T_40559;
  assign _GEN_5961 = {{16'd0}, _T_24454};
  assign _T_40599 = _GEN_5961 << 16;
  assign _GEN_5962 = {{8'd0}, _T_40563};
  assign _T_40603 = _GEN_5962 | _T_40599;
  assign _GEN_5963 = {{24'd0}, _T_24456};
  assign _T_40639 = _GEN_5963 << 24;
  assign _GEN_5964 = {{8'd0}, _T_40603};
  assign _T_40643 = _GEN_5964 | _T_40639;
  assign _GEN_5965 = {{8'd0}, _T_24556};
  assign _T_40719 = _GEN_5965 << 8;
  assign _GEN_5966 = {{8'd0}, _T_24554};
  assign _T_40723 = _GEN_5966 | _T_40719;
  assign _GEN_5967 = {{16'd0}, _T_24558};
  assign _T_40759 = _GEN_5967 << 16;
  assign _GEN_5968 = {{8'd0}, _T_40723};
  assign _T_40763 = _GEN_5968 | _T_40759;
  assign _GEN_5969 = {{24'd0}, _T_24560};
  assign _T_40799 = _GEN_5969 << 24;
  assign _GEN_5970 = {{8'd0}, _T_40763};
  assign _T_40803 = _GEN_5970 | _T_40799;
  assign _GEN_5971 = {{8'd0}, _T_25380};
  assign _T_40879 = _GEN_5971 << 8;
  assign _GEN_5972 = {{8'd0}, _T_25378};
  assign _T_40883 = _GEN_5972 | _T_40879;
  assign _GEN_5973 = {{16'd0}, _T_25382};
  assign _T_40919 = _GEN_5973 << 16;
  assign _GEN_5974 = {{8'd0}, _T_40883};
  assign _T_40923 = _GEN_5974 | _T_40919;
  assign _GEN_5975 = {{24'd0}, _T_25384};
  assign _T_40959 = _GEN_5975 << 24;
  assign _GEN_5976 = {{8'd0}, _T_40923};
  assign _T_40963 = _GEN_5976 | _T_40959;
  assign _GEN_5977 = {{8'd0}, _T_25068};
  assign _T_41039 = _GEN_5977 << 8;
  assign _GEN_5978 = {{8'd0}, _T_25066};
  assign _T_41043 = _GEN_5978 | _T_41039;
  assign _GEN_5979 = {{16'd0}, _T_25070};
  assign _T_41079 = _GEN_5979 << 16;
  assign _GEN_5980 = {{8'd0}, _T_41043};
  assign _T_41083 = _GEN_5980 | _T_41079;
  assign _GEN_5981 = {{24'd0}, _T_25072};
  assign _T_41119 = _GEN_5981 << 24;
  assign _GEN_5982 = {{8'd0}, _T_41083};
  assign _T_41123 = _GEN_5982 | _T_41119;
  assign _GEN_5983 = {{8'd0}, _T_23972};
  assign _T_41199 = _GEN_5983 << 8;
  assign _GEN_5984 = {{8'd0}, _T_23970};
  assign _T_41203 = _GEN_5984 | _T_41199;
  assign _GEN_5985 = {{16'd0}, _T_23974};
  assign _T_41239 = _GEN_5985 << 16;
  assign _GEN_5986 = {{8'd0}, _T_41203};
  assign _T_41243 = _GEN_5986 | _T_41239;
  assign _GEN_5987 = {{24'd0}, _T_23976};
  assign _T_41279 = _GEN_5987 << 24;
  assign _GEN_5988 = {{8'd0}, _T_41243};
  assign _T_41283 = _GEN_5988 | _T_41279;
  assign _GEN_5989 = {{8'd0}, _T_25028};
  assign _T_41359 = _GEN_5989 << 8;
  assign _GEN_5990 = {{8'd0}, _T_25026};
  assign _T_41363 = _GEN_5990 | _T_41359;
  assign _GEN_5991 = {{16'd0}, _T_25030};
  assign _T_41399 = _GEN_5991 << 16;
  assign _GEN_5992 = {{8'd0}, _T_41363};
  assign _T_41403 = _GEN_5992 | _T_41399;
  assign _GEN_5993 = {{24'd0}, _T_25032};
  assign _T_41439 = _GEN_5993 << 24;
  assign _GEN_5994 = {{8'd0}, _T_41403};
  assign _T_41443 = _GEN_5994 | _T_41439;
  assign _GEN_5995 = {{8'd0}, _T_24300};
  assign _T_41519 = _GEN_5995 << 8;
  assign _GEN_5996 = {{8'd0}, _T_24298};
  assign _T_41523 = _GEN_5996 | _T_41519;
  assign _GEN_5997 = {{16'd0}, _T_24302};
  assign _T_41559 = _GEN_5997 << 16;
  assign _GEN_5998 = {{8'd0}, _T_41523};
  assign _T_41563 = _GEN_5998 | _T_41559;
  assign _GEN_5999 = {{24'd0}, _T_24304};
  assign _T_41599 = _GEN_5999 << 24;
  assign _GEN_6000 = {{8'd0}, _T_41563};
  assign _T_41603 = _GEN_6000 | _T_41599;
  assign _GEN_6001 = {{8'd0}, _T_24012};
  assign _T_41679 = _GEN_6001 << 8;
  assign _GEN_6002 = {{8'd0}, _T_24010};
  assign _T_41683 = _GEN_6002 | _T_41679;
  assign _GEN_6003 = {{16'd0}, _T_24014};
  assign _T_41719 = _GEN_6003 << 16;
  assign _GEN_6004 = {{8'd0}, _T_41683};
  assign _T_41723 = _GEN_6004 | _T_41719;
  assign _GEN_6005 = {{24'd0}, _T_24016};
  assign _T_41759 = _GEN_6005 << 24;
  assign _GEN_6006 = {{8'd0}, _T_41723};
  assign _T_41763 = _GEN_6006 | _T_41759;
  assign _GEN_6007 = {{8'd0}, _T_25284};
  assign _T_41839 = _GEN_6007 << 8;
  assign _GEN_6008 = {{8'd0}, _T_25282};
  assign _T_41843 = _GEN_6008 | _T_41839;
  assign _GEN_6009 = {{16'd0}, _T_25286};
  assign _T_41879 = _GEN_6009 << 16;
  assign _GEN_6010 = {{8'd0}, _T_41843};
  assign _T_41883 = _GEN_6010 | _T_41879;
  assign _GEN_6011 = {{24'd0}, _T_25288};
  assign _T_41919 = _GEN_6011 << 24;
  assign _GEN_6012 = {{8'd0}, _T_41883};
  assign _T_41923 = _GEN_6012 | _T_41919;
  assign _GEN_6013 = {{8'd0}, _T_24228};
  assign _T_41999 = _GEN_6013 << 8;
  assign _GEN_6014 = {{8'd0}, _T_24226};
  assign _T_42003 = _GEN_6014 | _T_41999;
  assign _GEN_6015 = {{16'd0}, _T_24230};
  assign _T_42039 = _GEN_6015 << 16;
  assign _GEN_6016 = {{8'd0}, _T_42003};
  assign _T_42043 = _GEN_6016 | _T_42039;
  assign _GEN_6017 = {{24'd0}, _T_24232};
  assign _T_42079 = _GEN_6017 << 24;
  assign _GEN_6018 = {{8'd0}, _T_42043};
  assign _T_42083 = _GEN_6018 | _T_42079;
  assign _GEN_6019 = {{8'd0}, _T_23788};
  assign _T_42159 = _GEN_6019 << 8;
  assign _GEN_6020 = {{8'd0}, _T_23786};
  assign _T_42163 = _GEN_6020 | _T_42159;
  assign _GEN_6021 = {{16'd0}, _T_23790};
  assign _T_42199 = _GEN_6021 << 16;
  assign _GEN_6022 = {{8'd0}, _T_42163};
  assign _T_42203 = _GEN_6022 | _T_42199;
  assign _GEN_6023 = {{24'd0}, _T_23792};
  assign _T_42239 = _GEN_6023 << 24;
  assign _GEN_6024 = {{8'd0}, _T_42203};
  assign _T_42243 = _GEN_6024 | _T_42239;
  assign _T_42263 = _T_99490 & _T_35050;
  assign _GEN_2443 = _T_42263 ? _T_35064 : _GEN_353;
  assign _T_42303 = _T_99490 & _T_35090;
  assign _GEN_2444 = _T_42303 ? _T_35104 : _GEN_354;
  assign _T_42343 = _T_99490 & _T_35130;
  assign _GEN_2445 = _T_42343 ? _T_35144 : _GEN_355;
  assign _T_42383 = _T_99490 & _T_35170;
  assign _GEN_2446 = _T_42383 ? _T_35184 : _GEN_356;
  assign _GEN_6031 = {{8'd0}, _T_25500};
  assign _T_42479 = _GEN_6031 << 8;
  assign _GEN_6032 = {{8'd0}, _T_25498};
  assign _T_42483 = _GEN_6032 | _T_42479;
  assign _GEN_6033 = {{16'd0}, _T_25502};
  assign _T_42519 = _GEN_6033 << 16;
  assign _GEN_6034 = {{8'd0}, _T_42483};
  assign _T_42523 = _GEN_6034 | _T_42519;
  assign _GEN_6035 = {{24'd0}, _T_25504};
  assign _T_42559 = _GEN_6035 << 24;
  assign _GEN_6036 = {{8'd0}, _T_42523};
  assign _T_42563 = _GEN_6036 | _T_42559;
  assign _GEN_6037 = {{8'd0}, _T_25636};
  assign _T_42639 = _GEN_6037 << 8;
  assign _GEN_6038 = {{8'd0}, _T_25634};
  assign _T_42643 = _GEN_6038 | _T_42639;
  assign _GEN_6039 = {{16'd0}, _T_25638};
  assign _T_42679 = _GEN_6039 << 16;
  assign _GEN_6040 = {{8'd0}, _T_42643};
  assign _T_42683 = _GEN_6040 | _T_42679;
  assign _GEN_6041 = {{24'd0}, _T_25640};
  assign _T_42719 = _GEN_6041 << 24;
  assign _GEN_6042 = {{8'd0}, _T_42683};
  assign _T_42723 = _GEN_6042 | _T_42719;
  assign _GEN_6043 = {{8'd0}, _T_25244};
  assign _T_42799 = _GEN_6043 << 8;
  assign _GEN_6044 = {{8'd0}, _T_25242};
  assign _T_42803 = _GEN_6044 | _T_42799;
  assign _GEN_6045 = {{16'd0}, _T_25246};
  assign _T_42839 = _GEN_6045 << 16;
  assign _GEN_6046 = {{8'd0}, _T_42803};
  assign _T_42843 = _GEN_6046 | _T_42839;
  assign _GEN_6047 = {{24'd0}, _T_25248};
  assign _T_42879 = _GEN_6047 << 24;
  assign _GEN_6048 = {{8'd0}, _T_42843};
  assign _T_42883 = _GEN_6048 | _T_42879;
  assign _GEN_6049 = {{8'd0}, _T_24268};
  assign _T_42959 = _GEN_6049 << 8;
  assign _GEN_6050 = {{8'd0}, _T_24266};
  assign _T_42963 = _GEN_6050 | _T_42959;
  assign _GEN_6051 = {{16'd0}, _T_24270};
  assign _T_42999 = _GEN_6051 << 16;
  assign _GEN_6052 = {{8'd0}, _T_42963};
  assign _T_43003 = _GEN_6052 | _T_42999;
  assign _GEN_6053 = {{24'd0}, _T_24272};
  assign _T_43039 = _GEN_6053 << 24;
  assign _GEN_6054 = {{8'd0}, _T_43003};
  assign _T_43043 = _GEN_6054 | _T_43039;
  assign _GEN_6055 = {{8'd0}, _T_24708};
  assign _T_43119 = _GEN_6055 << 8;
  assign _GEN_6056 = {{8'd0}, _T_24706};
  assign _T_43123 = _GEN_6056 | _T_43119;
  assign _GEN_6057 = {{16'd0}, _T_24710};
  assign _T_43159 = _GEN_6057 << 16;
  assign _GEN_6058 = {{8'd0}, _T_43123};
  assign _T_43163 = _GEN_6058 | _T_43159;
  assign _GEN_6059 = {{24'd0}, _T_24712};
  assign _T_43199 = _GEN_6059 << 24;
  assign _GEN_6060 = {{8'd0}, _T_43163};
  assign _T_43203 = _GEN_6060 | _T_43199;
  assign _T_43223 = _T_99450 & _T_35050;
  assign _GEN_2447 = _T_43223 ? _T_35064 : _GEN_333;
  assign _T_43263 = _T_99450 & _T_35090;
  assign _GEN_2448 = _T_43263 ? _T_35104 : _GEN_334;
  assign _T_43303 = _T_99450 & _T_35130;
  assign _GEN_2449 = _T_43303 ? _T_35144 : _GEN_335;
  assign _T_43343 = _T_99450 & _T_35170;
  assign _GEN_2450 = _T_43343 ? _T_35184 : _GEN_336;
  assign _GEN_6067 = {{8'd0}, _T_25580};
  assign _T_43439 = _GEN_6067 << 8;
  assign _GEN_6068 = {{8'd0}, _T_25578};
  assign _T_43443 = _GEN_6068 | _T_43439;
  assign _GEN_6069 = {{16'd0}, _T_25582};
  assign _T_43479 = _GEN_6069 << 16;
  assign _GEN_6070 = {{8'd0}, _T_43443};
  assign _T_43483 = _GEN_6070 | _T_43479;
  assign _GEN_6071 = {{24'd0}, _T_25584};
  assign _T_43519 = _GEN_6071 << 24;
  assign _GEN_6072 = {{8'd0}, _T_43483};
  assign _T_43523 = _GEN_6072 | _T_43519;
  assign _GEN_6073 = {{8'd0}, _T_24484};
  assign _T_43759 = _GEN_6073 << 8;
  assign _GEN_6074 = {{8'd0}, _T_24482};
  assign _T_43763 = _GEN_6074 | _T_43759;
  assign _GEN_6075 = {{16'd0}, _T_24486};
  assign _T_43799 = _GEN_6075 << 16;
  assign _GEN_6076 = {{8'd0}, _T_43763};
  assign _T_43803 = _GEN_6076 | _T_43799;
  assign _GEN_6077 = {{24'd0}, _T_24488};
  assign _T_43839 = _GEN_6077 << 24;
  assign _GEN_6078 = {{8'd0}, _T_43803};
  assign _T_43843 = _GEN_6078 | _T_43839;
  assign _GEN_6079 = {{8'd0}, _T_24524};
  assign _T_43919 = _GEN_6079 << 8;
  assign _GEN_6080 = {{8'd0}, _T_24522};
  assign _T_43923 = _GEN_6080 | _T_43919;
  assign _GEN_6081 = {{16'd0}, _T_24526};
  assign _T_43959 = _GEN_6081 << 16;
  assign _GEN_6082 = {{8'd0}, _T_43923};
  assign _T_43963 = _GEN_6082 | _T_43959;
  assign _GEN_6083 = {{24'd0}, _T_24528};
  assign _T_43999 = _GEN_6083 << 24;
  assign _GEN_6084 = {{8'd0}, _T_43963};
  assign _T_44003 = _GEN_6084 | _T_43999;
  assign _GEN_6085 = {{8'd0}, _T_25540};
  assign _T_44079 = _GEN_6085 << 8;
  assign _GEN_6086 = {{8'd0}, _T_25538};
  assign _T_44083 = _GEN_6086 | _T_44079;
  assign _GEN_6087 = {{16'd0}, _T_25542};
  assign _T_44119 = _GEN_6087 << 16;
  assign _GEN_6088 = {{8'd0}, _T_44083};
  assign _T_44123 = _GEN_6088 | _T_44119;
  assign _GEN_6089 = {{24'd0}, _T_25544};
  assign _T_44159 = _GEN_6089 << 24;
  assign _GEN_6090 = {{8'd0}, _T_44123};
  assign _T_44163 = _GEN_6090 | _T_44159;
  assign _GEN_6091 = {{8'd0}, _T_24876};
  assign _T_44239 = _GEN_6091 << 8;
  assign _GEN_6092 = {{8'd0}, _T_24874};
  assign _T_44243 = _GEN_6092 | _T_44239;
  assign _GEN_6093 = {{16'd0}, _T_24878};
  assign _T_44279 = _GEN_6093 << 16;
  assign _GEN_6094 = {{8'd0}, _T_44243};
  assign _T_44283 = _GEN_6094 | _T_44279;
  assign _GEN_6095 = {{24'd0}, _T_24880};
  assign _T_44319 = _GEN_6095 << 24;
  assign _GEN_6096 = {{8'd0}, _T_44283};
  assign _T_44323 = _GEN_6096 | _T_44319;
  assign _GEN_6097 = {{8'd0}, _T_23940};
  assign _T_44399 = _GEN_6097 << 8;
  assign _GEN_6098 = {{8'd0}, _T_23938};
  assign _T_44403 = _GEN_6098 | _T_44399;
  assign _GEN_6099 = {{16'd0}, _T_23942};
  assign _T_44439 = _GEN_6099 << 16;
  assign _GEN_6100 = {{8'd0}, _T_44403};
  assign _T_44443 = _GEN_6100 | _T_44439;
  assign _GEN_6101 = {{24'd0}, _T_23944};
  assign _T_44479 = _GEN_6101 << 24;
  assign _GEN_6102 = {{8'd0}, _T_44443};
  assign _T_44483 = _GEN_6102 | _T_44479;
  assign _T_44503 = _T_99530 & _T_35050;
  assign _GEN_2451 = _T_44503 ? _T_35064 : _GEN_373;
  assign _T_44543 = _T_99530 & _T_35090;
  assign _GEN_2452 = _T_44543 ? _T_35104 : _GEN_374;
  assign _T_44583 = _T_99530 & _T_35130;
  assign _GEN_2453 = _T_44583 ? _T_35144 : _GEN_375;
  assign _T_44623 = _T_99530 & _T_35170;
  assign _GEN_2454 = _T_44623 ? _T_35184 : _GEN_376;
  assign _GEN_6109 = {{8'd0}, _T_24044};
  assign _T_44719 = _GEN_6109 << 8;
  assign _GEN_6110 = {{8'd0}, _T_24042};
  assign _T_44723 = _GEN_6110 | _T_44719;
  assign _GEN_6111 = {{16'd0}, _T_24046};
  assign _T_44759 = _GEN_6111 << 16;
  assign _GEN_6112 = {{8'd0}, _T_44723};
  assign _T_44763 = _GEN_6112 | _T_44759;
  assign _GEN_6113 = {{24'd0}, _T_24048};
  assign _T_44799 = _GEN_6113 << 24;
  assign _GEN_6114 = {{8'd0}, _T_44763};
  assign _T_44803 = _GEN_6114 | _T_44799;
  assign _GEN_6115 = {{8'd0}, _T_25324};
  assign _T_44879 = _GEN_6115 << 8;
  assign _GEN_6116 = {{8'd0}, _T_25322};
  assign _T_44883 = _GEN_6116 | _T_44879;
  assign _GEN_6117 = {{16'd0}, _T_25326};
  assign _T_44919 = _GEN_6117 << 16;
  assign _GEN_6118 = {{8'd0}, _T_44883};
  assign _T_44923 = _GEN_6118 | _T_44919;
  assign _GEN_6119 = {{24'd0}, _T_25328};
  assign _T_44959 = _GEN_6119 << 24;
  assign _GEN_6120 = {{8'd0}, _T_44923};
  assign _T_44963 = _GEN_6120 | _T_44959;
  assign _GEN_6121 = {{8'd0}, _T_24868};
  assign _T_45039 = _GEN_6121 << 8;
  assign _GEN_6122 = {{8'd0}, _T_24866};
  assign _T_45043 = _GEN_6122 | _T_45039;
  assign _GEN_6123 = {{16'd0}, _T_24870};
  assign _T_45079 = _GEN_6123 << 16;
  assign _GEN_6124 = {{8'd0}, _T_45043};
  assign _T_45083 = _GEN_6124 | _T_45079;
  assign _GEN_6125 = {{24'd0}, _T_24872};
  assign _T_45119 = _GEN_6125 << 24;
  assign _GEN_6126 = {{8'd0}, _T_45083};
  assign _T_45123 = _GEN_6126 | _T_45119;
  assign _GEN_6127 = {{8'd0}, _T_24988};
  assign _T_45199 = _GEN_6127 << 8;
  assign _GEN_6128 = {{8'd0}, _T_24986};
  assign _T_45203 = _GEN_6128 | _T_45199;
  assign _GEN_6129 = {{16'd0}, _T_24990};
  assign _T_45239 = _GEN_6129 << 16;
  assign _GEN_6130 = {{8'd0}, _T_45203};
  assign _T_45243 = _GEN_6130 | _T_45239;
  assign _GEN_6131 = {{24'd0}, _T_24992};
  assign _T_45279 = _GEN_6131 << 24;
  assign _GEN_6132 = {{8'd0}, _T_45243};
  assign _T_45283 = _GEN_6132 | _T_45279;
  assign _GEN_6133 = {{8'd0}, _T_25124};
  assign _T_45359 = _GEN_6133 << 8;
  assign _GEN_6134 = {{8'd0}, _T_25122};
  assign _T_45363 = _GEN_6134 | _T_45359;
  assign _GEN_6135 = {{16'd0}, _T_25126};
  assign _T_45399 = _GEN_6135 << 16;
  assign _GEN_6136 = {{8'd0}, _T_45363};
  assign _T_45403 = _GEN_6136 | _T_45399;
  assign _GEN_6137 = {{24'd0}, _T_25128};
  assign _T_45439 = _GEN_6137 << 24;
  assign _GEN_6138 = {{8'd0}, _T_45403};
  assign _T_45443 = _GEN_6138 | _T_45439;
  assign _GEN_6139 = {{8'd0}, _T_23820};
  assign _T_45519 = _GEN_6139 << 8;
  assign _GEN_6140 = {{8'd0}, _T_23818};
  assign _T_45523 = _GEN_6140 | _T_45519;
  assign _GEN_6141 = {{16'd0}, _T_23822};
  assign _T_45559 = _GEN_6141 << 16;
  assign _GEN_6142 = {{8'd0}, _T_45523};
  assign _T_45563 = _GEN_6142 | _T_45559;
  assign _GEN_6143 = {{24'd0}, _T_23824};
  assign _T_45599 = _GEN_6143 << 24;
  assign _GEN_6144 = {{8'd0}, _T_45563};
  assign _T_45603 = _GEN_6144 | _T_45599;
  assign _GEN_6145 = {{8'd0}, _T_25756};
  assign _T_45679 = _GEN_6145 << 8;
  assign _GEN_6146 = {{8'd0}, _T_25754};
  assign _T_45683 = _GEN_6146 | _T_45679;
  assign _GEN_6147 = {{16'd0}, _T_25758};
  assign _T_45719 = _GEN_6147 << 16;
  assign _GEN_6148 = {{8'd0}, _T_45683};
  assign _T_45723 = _GEN_6148 | _T_45719;
  assign _GEN_6149 = {{24'd0}, _T_25760};
  assign _T_45759 = _GEN_6149 << 24;
  assign _GEN_6150 = {{8'd0}, _T_45723};
  assign _T_45763 = _GEN_6150 | _T_45759;
  assign _GEN_6151 = {{8'd0}, _T_24196};
  assign _T_45999 = _GEN_6151 << 8;
  assign _GEN_6152 = {{8'd0}, _T_24194};
  assign _T_46003 = _GEN_6152 | _T_45999;
  assign _GEN_6153 = {{16'd0}, _T_24198};
  assign _T_46039 = _GEN_6153 << 16;
  assign _GEN_6154 = {{8'd0}, _T_46003};
  assign _T_46043 = _GEN_6154 | _T_46039;
  assign _GEN_6155 = {{24'd0}, _T_24200};
  assign _T_46079 = _GEN_6155 << 24;
  assign _GEN_6156 = {{8'd0}, _T_46043};
  assign _T_46083 = _GEN_6156 | _T_46079;
  assign _GEN_6157 = {{8'd0}, _T_24156};
  assign _T_46199 = _GEN_6157 << 8;
  assign _GEN_6158 = {{8'd0}, _T_24154};
  assign _T_46203 = _GEN_6158 | _T_46199;
  assign _GEN_6159 = {{16'd0}, _T_24158};
  assign _T_46239 = _GEN_6159 << 16;
  assign _GEN_6160 = {{8'd0}, _T_46203};
  assign _T_46243 = _GEN_6160 | _T_46239;
  assign _GEN_6161 = {{24'd0}, _T_24160};
  assign _T_46279 = _GEN_6161 << 24;
  assign _GEN_6162 = {{8'd0}, _T_46243};
  assign _T_46283 = _GEN_6162 | _T_46279;
  assign _GEN_6163 = {{8'd0}, _T_24036};
  assign _T_46359 = _GEN_6163 << 8;
  assign _GEN_6164 = {{8'd0}, _T_24034};
  assign _T_46363 = _GEN_6164 | _T_46359;
  assign _GEN_6165 = {{16'd0}, _T_24038};
  assign _T_46399 = _GEN_6165 << 16;
  assign _GEN_6166 = {{8'd0}, _T_46363};
  assign _T_46403 = _GEN_6166 | _T_46399;
  assign _GEN_6167 = {{24'd0}, _T_24040};
  assign _T_46439 = _GEN_6167 << 24;
  assign _GEN_6168 = {{8'd0}, _T_46403};
  assign _T_46443 = _GEN_6168 | _T_46439;
  assign _GEN_6169 = {{8'd0}, _T_25316};
  assign _T_46519 = _GEN_6169 << 8;
  assign _GEN_6170 = {{8'd0}, _T_25314};
  assign _T_46523 = _GEN_6170 | _T_46519;
  assign _GEN_6171 = {{16'd0}, _T_25318};
  assign _T_46559 = _GEN_6171 << 16;
  assign _GEN_6172 = {{8'd0}, _T_46523};
  assign _T_46563 = _GEN_6172 | _T_46559;
  assign _GEN_6173 = {{24'd0}, _T_25320};
  assign _T_46599 = _GEN_6173 << 24;
  assign _GEN_6174 = {{8'd0}, _T_46563};
  assign _T_46603 = _GEN_6174 | _T_46599;
  assign _GEN_6175 = {{8'd0}, _T_24740};
  assign _T_46679 = _GEN_6175 << 8;
  assign _GEN_6176 = {{8'd0}, _T_24738};
  assign _T_46683 = _GEN_6176 | _T_46679;
  assign _GEN_6177 = {{16'd0}, _T_24742};
  assign _T_46719 = _GEN_6177 << 16;
  assign _GEN_6178 = {{8'd0}, _T_46683};
  assign _T_46723 = _GEN_6178 | _T_46719;
  assign _GEN_6179 = {{24'd0}, _T_24744};
  assign _T_46759 = _GEN_6179 << 24;
  assign _GEN_6180 = {{8'd0}, _T_46723};
  assign _T_46763 = _GEN_6180 | _T_46759;
  assign _GEN_6181 = {{8'd0}, _T_25212};
  assign _T_46999 = _GEN_6181 << 8;
  assign _GEN_6182 = {{8'd0}, _T_25210};
  assign _T_47003 = _GEN_6182 | _T_46999;
  assign _GEN_6183 = {{16'd0}, _T_25214};
  assign _T_47039 = _GEN_6183 << 16;
  assign _GEN_6184 = {{8'd0}, _T_47003};
  assign _T_47043 = _GEN_6184 | _T_47039;
  assign _GEN_6185 = {{24'd0}, _T_25216};
  assign _T_47079 = _GEN_6185 << 24;
  assign _GEN_6186 = {{8'd0}, _T_47043};
  assign _T_47083 = _GEN_6186 | _T_47079;
  assign _GEN_6187 = {{8'd0}, _T_23860};
  assign _T_47159 = _GEN_6187 << 8;
  assign _GEN_6188 = {{8'd0}, _T_23858};
  assign _T_47163 = _GEN_6188 | _T_47159;
  assign _GEN_6189 = {{16'd0}, _T_23862};
  assign _T_47199 = _GEN_6189 << 16;
  assign _GEN_6190 = {{8'd0}, _T_47163};
  assign _T_47203 = _GEN_6190 | _T_47199;
  assign _GEN_6191 = {{24'd0}, _T_23864};
  assign _T_47239 = _GEN_6191 << 24;
  assign _GEN_6192 = {{8'd0}, _T_47203};
  assign _T_47243 = _GEN_6192 | _T_47239;
  assign _GEN_6193 = {{8'd0}, _T_24748};
  assign _T_47479 = _GEN_6193 << 8;
  assign _GEN_6194 = {{8'd0}, _T_24746};
  assign _T_47483 = _GEN_6194 | _T_47479;
  assign _GEN_6195 = {{16'd0}, _T_24750};
  assign _T_47519 = _GEN_6195 << 16;
  assign _GEN_6196 = {{8'd0}, _T_47483};
  assign _T_47523 = _GEN_6196 | _T_47519;
  assign _GEN_6197 = {{24'd0}, _T_24752};
  assign _T_47559 = _GEN_6197 << 24;
  assign _GEN_6198 = {{8'd0}, _T_47523};
  assign _T_47563 = _GEN_6198 | _T_47559;
  assign _T_47583 = _T_99522 & _T_35050;
  assign _GEN_2455 = _T_47583 ? _T_35064 : _GEN_369;
  assign _T_47623 = _T_99522 & _T_35090;
  assign _GEN_2456 = _T_47623 ? _T_35104 : _GEN_370;
  assign _T_47663 = _T_99522 & _T_35130;
  assign _GEN_2457 = _T_47663 ? _T_35144 : _GEN_371;
  assign _T_47703 = _T_99522 & _T_35170;
  assign _GEN_2458 = _T_47703 ? _T_35184 : _GEN_372;
  assign _GEN_6205 = {{8'd0}, _T_24628};
  assign _T_47799 = _GEN_6205 << 8;
  assign _GEN_6206 = {{8'd0}, _T_24626};
  assign _T_47803 = _GEN_6206 | _T_47799;
  assign _GEN_6207 = {{16'd0}, _T_24630};
  assign _T_47839 = _GEN_6207 << 16;
  assign _GEN_6208 = {{8'd0}, _T_47803};
  assign _T_47843 = _GEN_6208 | _T_47839;
  assign _GEN_6209 = {{24'd0}, _T_24632};
  assign _T_47879 = _GEN_6209 << 24;
  assign _GEN_6210 = {{8'd0}, _T_47843};
  assign _T_47883 = _GEN_6210 | _T_47879;
  assign _GEN_6211 = {{8'd0}, _T_24372};
  assign _T_48119 = _GEN_6211 << 8;
  assign _GEN_6212 = {{8'd0}, _T_24370};
  assign _T_48123 = _GEN_6212 | _T_48119;
  assign _GEN_6213 = {{16'd0}, _T_24374};
  assign _T_48159 = _GEN_6213 << 16;
  assign _GEN_6214 = {{8'd0}, _T_48123};
  assign _T_48163 = _GEN_6214 | _T_48159;
  assign _GEN_6215 = {{24'd0}, _T_24376};
  assign _T_48199 = _GEN_6215 << 24;
  assign _GEN_6216 = {{8'd0}, _T_48163};
  assign _T_48203 = _GEN_6216 | _T_48199;
  assign _GEN_6217 = {{8'd0}, _T_24116};
  assign _T_48279 = _GEN_6217 << 8;
  assign _GEN_6218 = {{8'd0}, _T_24114};
  assign _T_48283 = _GEN_6218 | _T_48279;
  assign _GEN_6219 = {{16'd0}, _T_24118};
  assign _T_48319 = _GEN_6219 << 16;
  assign _GEN_6220 = {{8'd0}, _T_48283};
  assign _T_48323 = _GEN_6220 | _T_48319;
  assign _GEN_6221 = {{24'd0}, _T_24120};
  assign _T_48359 = _GEN_6221 << 24;
  assign _GEN_6222 = {{8'd0}, _T_48323};
  assign _T_48363 = _GEN_6222 | _T_48359;
  assign _GEN_6223 = {{8'd0}, _T_23780};
  assign _T_48439 = _GEN_6223 << 8;
  assign _GEN_6224 = {{8'd0}, _T_23778};
  assign _T_48443 = _GEN_6224 | _T_48439;
  assign _GEN_6225 = {{16'd0}, _T_23782};
  assign _T_48479 = _GEN_6225 << 16;
  assign _GEN_6226 = {{8'd0}, _T_48443};
  assign _T_48483 = _GEN_6226 | _T_48479;
  assign _GEN_6227 = {{24'd0}, _T_23784};
  assign _T_48519 = _GEN_6227 << 24;
  assign _GEN_6228 = {{8'd0}, _T_48483};
  assign _T_48523 = _GEN_6228 | _T_48519;
  assign _GEN_6229 = {{8'd0}, _T_24492};
  assign _T_48599 = _GEN_6229 << 8;
  assign _GEN_6230 = {{8'd0}, _T_24490};
  assign _T_48603 = _GEN_6230 | _T_48599;
  assign _GEN_6231 = {{16'd0}, _T_24494};
  assign _T_48639 = _GEN_6231 << 16;
  assign _GEN_6232 = {{8'd0}, _T_48603};
  assign _T_48643 = _GEN_6232 | _T_48639;
  assign _GEN_6233 = {{24'd0}, _T_24496};
  assign _T_48679 = _GEN_6233 << 24;
  assign _GEN_6234 = {{8'd0}, _T_48643};
  assign _T_48683 = _GEN_6234 | _T_48679;
  assign _GEN_6235 = {{8'd0}, _T_24836};
  assign _T_48759 = _GEN_6235 << 8;
  assign _GEN_6236 = {{8'd0}, _T_24834};
  assign _T_48763 = _GEN_6236 | _T_48759;
  assign _GEN_6237 = {{16'd0}, _T_24838};
  assign _T_48799 = _GEN_6237 << 16;
  assign _GEN_6238 = {{8'd0}, _T_48763};
  assign _T_48803 = _GEN_6238 | _T_48799;
  assign _GEN_6239 = {{24'd0}, _T_24840};
  assign _T_48839 = _GEN_6239 << 24;
  assign _GEN_6240 = {{8'd0}, _T_48803};
  assign _T_48843 = _GEN_6240 | _T_48839;
  assign _GEN_6241 = {{8'd0}, _T_24076};
  assign _T_48919 = _GEN_6241 << 8;
  assign _GEN_6242 = {{8'd0}, _T_24074};
  assign _T_48923 = _GEN_6242 | _T_48919;
  assign _GEN_6243 = {{16'd0}, _T_24078};
  assign _T_48959 = _GEN_6243 << 16;
  assign _GEN_6244 = {{8'd0}, _T_48923};
  assign _T_48963 = _GEN_6244 | _T_48959;
  assign _GEN_6245 = {{24'd0}, _T_24080};
  assign _T_48999 = _GEN_6245 << 24;
  assign _GEN_6246 = {{8'd0}, _T_48963};
  assign _T_49003 = _GEN_6246 | _T_48999;
  assign _GEN_6247 = {{8'd0}, _T_25092};
  assign _T_49079 = _GEN_6247 << 8;
  assign _GEN_6248 = {{8'd0}, _T_25090};
  assign _T_49083 = _GEN_6248 | _T_49079;
  assign _GEN_6249 = {{16'd0}, _T_25094};
  assign _T_49119 = _GEN_6249 << 16;
  assign _GEN_6250 = {{8'd0}, _T_49083};
  assign _T_49123 = _GEN_6250 | _T_49119;
  assign _GEN_6251 = {{24'd0}, _T_25096};
  assign _T_49159 = _GEN_6251 << 24;
  assign _GEN_6252 = {{8'd0}, _T_49123};
  assign _T_49163 = _GEN_6252 | _T_49159;
  assign _GEN_6253 = {{8'd0}, _T_24956};
  assign _T_49279 = _GEN_6253 << 8;
  assign _GEN_6254 = {{8'd0}, _T_24954};
  assign _T_49283 = _GEN_6254 | _T_49279;
  assign _GEN_6255 = {{16'd0}, _T_24958};
  assign _T_49319 = _GEN_6255 << 16;
  assign _GEN_6256 = {{8'd0}, _T_49283};
  assign _T_49323 = _GEN_6256 | _T_49319;
  assign _GEN_6257 = {{24'd0}, _T_24960};
  assign _T_49359 = _GEN_6257 << 24;
  assign _GEN_6258 = {{8'd0}, _T_49323};
  assign _T_49363 = _GEN_6258 | _T_49359;
  assign _GEN_6259 = {{8'd0}, _T_25132};
  assign _T_49439 = _GEN_6259 << 8;
  assign _GEN_6260 = {{8'd0}, _T_25130};
  assign _T_49443 = _GEN_6260 | _T_49439;
  assign _GEN_6261 = {{16'd0}, _T_25134};
  assign _T_49479 = _GEN_6261 << 16;
  assign _GEN_6262 = {{8'd0}, _T_49443};
  assign _T_49483 = _GEN_6262 | _T_49479;
  assign _GEN_6263 = {{24'd0}, _T_25136};
  assign _T_49519 = _GEN_6263 << 24;
  assign _GEN_6264 = {{8'd0}, _T_49483};
  assign _T_49523 = _GEN_6264 | _T_49519;
  assign _GEN_6265 = {{8'd0}, _T_23900};
  assign _T_49599 = _GEN_6265 << 8;
  assign _GEN_6266 = {{8'd0}, _T_23898};
  assign _T_49603 = _GEN_6266 | _T_49599;
  assign _GEN_6267 = {{16'd0}, _T_23902};
  assign _T_49639 = _GEN_6267 << 16;
  assign _GEN_6268 = {{8'd0}, _T_49603};
  assign _T_49643 = _GEN_6268 | _T_49639;
  assign _GEN_6269 = {{24'd0}, _T_23904};
  assign _T_49679 = _GEN_6269 << 24;
  assign _GEN_6270 = {{8'd0}, _T_49643};
  assign _T_49683 = _GEN_6270 | _T_49679;
  assign _GEN_6271 = {{8'd0}, _T_25436};
  assign _T_49759 = _GEN_6271 << 8;
  assign _GEN_6272 = {{8'd0}, _T_25434};
  assign _T_49763 = _GEN_6272 | _T_49759;
  assign _GEN_6273 = {{16'd0}, _T_25438};
  assign _T_49799 = _GEN_6273 << 16;
  assign _GEN_6274 = {{8'd0}, _T_49763};
  assign _T_49803 = _GEN_6274 | _T_49799;
  assign _GEN_6275 = {{24'd0}, _T_25440};
  assign _T_49839 = _GEN_6275 << 24;
  assign _GEN_6276 = {{8'd0}, _T_49803};
  assign _T_49843 = _GEN_6276 | _T_49839;
  assign _GEN_6277 = {{8'd0}, _T_25572};
  assign _T_49919 = _GEN_6277 << 8;
  assign _GEN_6278 = {{8'd0}, _T_25570};
  assign _T_49923 = _GEN_6278 | _T_49919;
  assign _GEN_6279 = {{16'd0}, _T_25574};
  assign _T_49959 = _GEN_6279 << 16;
  assign _GEN_6280 = {{8'd0}, _T_49923};
  assign _T_49963 = _GEN_6280 | _T_49959;
  assign _GEN_6281 = {{24'd0}, _T_25576};
  assign _T_49999 = _GEN_6281 << 24;
  assign _GEN_6282 = {{8'd0}, _T_49963};
  assign _T_50003 = _GEN_6282 | _T_49999;
  assign _GEN_6283 = {{8'd0}, _T_24588};
  assign _T_50079 = _GEN_6283 << 8;
  assign _GEN_6284 = {{8'd0}, _T_24586};
  assign _T_50083 = _GEN_6284 | _T_50079;
  assign _GEN_6285 = {{16'd0}, _T_24590};
  assign _T_50119 = _GEN_6285 << 16;
  assign _GEN_6286 = {{8'd0}, _T_50083};
  assign _T_50123 = _GEN_6286 | _T_50119;
  assign _GEN_6287 = {{24'd0}, _T_24592};
  assign _T_50159 = _GEN_6287 << 24;
  assign _GEN_6288 = {{8'd0}, _T_50123};
  assign _T_50163 = _GEN_6288 | _T_50159;
  assign _T_50164 = _T_35020[9:0];
  assign _T_50168 = ~ _T_50164;
  assign _T_50170 = _T_50168 == 10'h0;
  assign _T_50183 = _T_98282 & _T_50170;
  assign _T_50184 = io_hart_in_0_a_bits_data[9:0];
  assign _GEN_6289 = {{8'd0}, _T_25180};
  assign _T_50279 = _GEN_6289 << 8;
  assign _GEN_6290 = {{8'd0}, _T_25178};
  assign _T_50283 = _GEN_6290 | _T_50279;
  assign _GEN_6291 = {{16'd0}, _T_25182};
  assign _T_50319 = _GEN_6291 << 16;
  assign _GEN_6292 = {{8'd0}, _T_50283};
  assign _T_50323 = _GEN_6292 | _T_50319;
  assign _GEN_6293 = {{24'd0}, _T_25184};
  assign _T_50359 = _GEN_6293 << 24;
  assign _GEN_6294 = {{8'd0}, _T_50323};
  assign _T_50363 = _GEN_6294 | _T_50359;
  assign _GEN_6295 = {{8'd0}, _T_24332};
  assign _T_50439 = _GEN_6295 << 8;
  assign _GEN_6296 = {{8'd0}, _T_24330};
  assign _T_50443 = _GEN_6296 | _T_50439;
  assign _GEN_6297 = {{16'd0}, _T_24334};
  assign _T_50479 = _GEN_6297 << 16;
  assign _GEN_6298 = {{8'd0}, _T_50443};
  assign _T_50483 = _GEN_6298 | _T_50479;
  assign _GEN_6299 = {{24'd0}, _T_24336};
  assign _T_50519 = _GEN_6299 << 24;
  assign _GEN_6300 = {{8'd0}, _T_50483};
  assign _T_50523 = _GEN_6300 | _T_50519;
  assign _GEN_6301 = {{8'd0}, _T_25388};
  assign _T_50759 = _GEN_6301 << 8;
  assign _GEN_6302 = {{8'd0}, _T_25386};
  assign _T_50763 = _GEN_6302 | _T_50759;
  assign _GEN_6303 = {{16'd0}, _T_25390};
  assign _T_50799 = _GEN_6303 << 16;
  assign _GEN_6304 = {{8'd0}, _T_50763};
  assign _T_50803 = _GEN_6304 | _T_50799;
  assign _GEN_6305 = {{24'd0}, _T_25392};
  assign _T_50839 = _GEN_6305 << 24;
  assign _GEN_6306 = {{8'd0}, _T_50803};
  assign _T_50843 = _GEN_6306 | _T_50839;
  assign _GEN_6307 = {{8'd0}, _T_25644};
  assign _T_50919 = _GEN_6307 << 8;
  assign _GEN_6308 = {{8'd0}, _T_25642};
  assign _T_50923 = _GEN_6308 | _T_50919;
  assign _GEN_6309 = {{16'd0}, _T_25646};
  assign _T_50959 = _GEN_6309 << 16;
  assign _GEN_6310 = {{8'd0}, _T_50923};
  assign _T_50963 = _GEN_6310 | _T_50959;
  assign _GEN_6311 = {{24'd0}, _T_25648};
  assign _T_50999 = _GEN_6311 << 24;
  assign _GEN_6312 = {{8'd0}, _T_50963};
  assign _T_51003 = _GEN_6312 | _T_50999;
  assign _GEN_6313 = {{8'd0}, _T_25348};
  assign _T_51079 = _GEN_6313 << 8;
  assign _GEN_6314 = {{8'd0}, _T_25346};
  assign _T_51083 = _GEN_6314 | _T_51079;
  assign _GEN_6315 = {{16'd0}, _T_25350};
  assign _T_51119 = _GEN_6315 << 16;
  assign _GEN_6316 = {{8'd0}, _T_51083};
  assign _T_51123 = _GEN_6316 | _T_51119;
  assign _GEN_6317 = {{24'd0}, _T_25352};
  assign _T_51159 = _GEN_6317 << 24;
  assign _GEN_6318 = {{8'd0}, _T_51123};
  assign _T_51163 = _GEN_6318 | _T_51159;
  assign _GEN_6319 = {{8'd0}, _T_24292};
  assign _T_51239 = _GEN_6319 << 8;
  assign _GEN_6320 = {{8'd0}, _T_24290};
  assign _T_51243 = _GEN_6320 | _T_51239;
  assign _GEN_6321 = {{16'd0}, _T_24294};
  assign _T_51279 = _GEN_6321 << 16;
  assign _GEN_6322 = {{8'd0}, _T_51243};
  assign _T_51283 = _GEN_6322 | _T_51279;
  assign _GEN_6323 = {{24'd0}, _T_24296};
  assign _T_51319 = _GEN_6323 << 24;
  assign _GEN_6324 = {{8'd0}, _T_51283};
  assign _T_51323 = _GEN_6324 | _T_51319;
  assign _GEN_6325 = {{8'd0}, _T_23980};
  assign _T_51399 = _GEN_6325 << 8;
  assign _GEN_6326 = {{8'd0}, _T_23978};
  assign _T_51403 = _GEN_6326 | _T_51399;
  assign _GEN_6327 = {{16'd0}, _T_23982};
  assign _T_51439 = _GEN_6327 << 16;
  assign _GEN_6328 = {{8'd0}, _T_51403};
  assign _T_51443 = _GEN_6328 | _T_51439;
  assign _GEN_6329 = {{24'd0}, _T_23984};
  assign _T_51479 = _GEN_6329 << 24;
  assign _GEN_6330 = {{8'd0}, _T_51443};
  assign _T_51483 = _GEN_6330 | _T_51479;
  assign _T_51503 = _T_99554 & _T_35050;
  assign _GEN_2460 = _T_51503 ? _T_35064 : _GEN_317;
  assign _T_51543 = _T_99554 & _T_35090;
  assign _GEN_2461 = _T_51543 ? _T_35104 : _GEN_318;
  assign _T_51583 = _T_99554 & _T_35130;
  assign _GEN_2462 = _T_51583 ? _T_35144 : _GEN_319;
  assign _T_51623 = _T_99554 & _T_35170;
  assign _GEN_2463 = _T_51623 ? _T_35184 : _GEN_320;
  assign _GEN_6337 = {{8'd0}, _T_24236};
  assign _T_51879 = _GEN_6337 << 8;
  assign _GEN_6338 = {{8'd0}, _T_24234};
  assign _T_51883 = _GEN_6338 | _T_51879;
  assign _GEN_6339 = {{16'd0}, _T_24238};
  assign _T_51919 = _GEN_6339 << 16;
  assign _GEN_6340 = {{8'd0}, _T_51883};
  assign _T_51923 = _GEN_6340 | _T_51919;
  assign _GEN_6341 = {{24'd0}, _T_24240};
  assign _T_51959 = _GEN_6341 << 24;
  assign _GEN_6342 = {{8'd0}, _T_51923};
  assign _T_51963 = _GEN_6342 | _T_51959;
  assign _GEN_6343 = {{8'd0}, _T_24924};
  assign _T_52039 = _GEN_6343 << 8;
  assign _GEN_6344 = {{8'd0}, _T_24922};
  assign _T_52043 = _GEN_6344 | _T_52039;
  assign _GEN_6345 = {{16'd0}, _T_24926};
  assign _T_52079 = _GEN_6345 << 16;
  assign _GEN_6346 = {{8'd0}, _T_52043};
  assign _T_52083 = _GEN_6346 | _T_52079;
  assign _GEN_6347 = {{24'd0}, _T_24928};
  assign _T_52119 = _GEN_6347 << 24;
  assign _GEN_6348 = {{8'd0}, _T_52083};
  assign _T_52123 = _GEN_6348 | _T_52119;
  assign _GEN_6349 = {{8'd0}, _T_24804};
  assign _T_52199 = _GEN_6349 << 8;
  assign _GEN_6350 = {{8'd0}, _T_24802};
  assign _T_52203 = _GEN_6350 | _T_52199;
  assign _GEN_6351 = {{16'd0}, _T_24806};
  assign _T_52239 = _GEN_6351 << 16;
  assign _GEN_6352 = {{8'd0}, _T_52203};
  assign _T_52243 = _GEN_6352 | _T_52239;
  assign _GEN_6353 = {{24'd0}, _T_24808};
  assign _T_52279 = _GEN_6353 << 24;
  assign _GEN_6354 = {{8'd0}, _T_52243};
  assign _T_52283 = _GEN_6354 | _T_52279;
  assign _GEN_6355 = {{8'd0}, _T_24548};
  assign _T_52359 = _GEN_6355 << 8;
  assign _GEN_6356 = {{8'd0}, _T_24546};
  assign _T_52363 = _GEN_6356 | _T_52359;
  assign _GEN_6357 = {{16'd0}, _T_24550};
  assign _T_52399 = _GEN_6357 << 16;
  assign _GEN_6358 = {{8'd0}, _T_52363};
  assign _T_52403 = _GEN_6358 | _T_52399;
  assign _GEN_6359 = {{24'd0}, _T_24552};
  assign _T_52439 = _GEN_6359 << 24;
  assign _GEN_6360 = {{8'd0}, _T_52403};
  assign _T_52443 = _GEN_6360 | _T_52439;
  assign _GEN_6361 = {{8'd0}, _T_25060};
  assign _T_52519 = _GEN_6361 << 8;
  assign _GEN_6362 = {{8'd0}, _T_25058};
  assign _T_52523 = _GEN_6362 | _T_52519;
  assign _GEN_6363 = {{16'd0}, _T_25062};
  assign _T_52559 = _GEN_6363 << 16;
  assign _GEN_6364 = {{8'd0}, _T_52523};
  assign _T_52563 = _GEN_6364 | _T_52559;
  assign _GEN_6365 = {{24'd0}, _T_25064};
  assign _T_52599 = _GEN_6365 << 24;
  assign _GEN_6366 = {{8'd0}, _T_52563};
  assign _T_52603 = _GEN_6366 | _T_52599;
  assign _GEN_6367 = {{8'd0}, _T_25692};
  assign _T_52679 = _GEN_6367 << 8;
  assign _GEN_6368 = {{8'd0}, _T_25690};
  assign _T_52683 = _GEN_6368 | _T_52679;
  assign _GEN_6369 = {{16'd0}, _T_25694};
  assign _T_52719 = _GEN_6369 << 16;
  assign _GEN_6370 = {{8'd0}, _T_52683};
  assign _T_52723 = _GEN_6370 | _T_52719;
  assign _GEN_6371 = {{24'd0}, _T_25696};
  assign _T_52759 = _GEN_6371 << 24;
  assign _GEN_6372 = {{8'd0}, _T_52723};
  assign _T_52763 = _GEN_6372 | _T_52759;
  assign _GEN_6373 = {{8'd0}, _T_24324};
  assign _T_52839 = _GEN_6373 << 8;
  assign _GEN_6374 = {{8'd0}, _T_24322};
  assign _T_52843 = _GEN_6374 | _T_52839;
  assign _GEN_6375 = {{16'd0}, _T_24326};
  assign _T_52879 = _GEN_6375 << 16;
  assign _GEN_6376 = {{8'd0}, _T_52843};
  assign _T_52883 = _GEN_6376 | _T_52879;
  assign _GEN_6377 = {{24'd0}, _T_24328};
  assign _T_52919 = _GEN_6377 << 24;
  assign _GEN_6378 = {{8'd0}, _T_52883};
  assign _T_52923 = _GEN_6378 | _T_52919;
  assign _GEN_6379 = {{8'd0}, _T_25468};
  assign _T_52999 = _GEN_6379 << 8;
  assign _GEN_6380 = {{8'd0}, _T_25466};
  assign _T_53003 = _GEN_6380 | _T_52999;
  assign _GEN_6381 = {{16'd0}, _T_25470};
  assign _T_53039 = _GEN_6381 << 16;
  assign _GEN_6382 = {{8'd0}, _T_53003};
  assign _T_53043 = _GEN_6382 | _T_53039;
  assign _GEN_6383 = {{24'd0}, _T_25472};
  assign _T_53079 = _GEN_6383 << 24;
  assign _GEN_6384 = {{8'd0}, _T_53043};
  assign _T_53083 = _GEN_6384 | _T_53079;
  assign _GEN_6385 = {{8'd0}, _T_23748};
  assign _T_53159 = _GEN_6385 << 8;
  assign _GEN_6386 = {{8'd0}, _T_23746};
  assign _T_53163 = _GEN_6386 | _T_53159;
  assign _GEN_6387 = {{16'd0}, _T_23750};
  assign _T_53199 = _GEN_6387 << 16;
  assign _GEN_6388 = {{8'd0}, _T_53163};
  assign _T_53203 = _GEN_6388 | _T_53199;
  assign _GEN_6389 = {{24'd0}, _T_23752};
  assign _T_53239 = _GEN_6389 << 24;
  assign _GEN_6390 = {{8'd0}, _T_53203};
  assign _T_53243 = _GEN_6390 | _T_53239;
  assign _GEN_6391 = {{8'd0}, _T_25604};
  assign _T_53319 = _GEN_6391 << 8;
  assign _GEN_6392 = {{8'd0}, _T_25602};
  assign _T_53323 = _GEN_6392 | _T_53319;
  assign _GEN_6393 = {{16'd0}, _T_25606};
  assign _T_53359 = _GEN_6393 << 16;
  assign _GEN_6394 = {{8'd0}, _T_53323};
  assign _T_53363 = _GEN_6394 | _T_53359;
  assign _GEN_6395 = {{24'd0}, _T_25608};
  assign _T_53399 = _GEN_6395 << 24;
  assign _GEN_6396 = {{8'd0}, _T_53363};
  assign _T_53403 = _GEN_6396 | _T_53399;
  assign _GEN_6397 = {{8'd0}, _T_24412};
  assign _T_53479 = _GEN_6397 << 8;
  assign _GEN_6398 = {{8'd0}, _T_24410};
  assign _T_53483 = _GEN_6398 | _T_53479;
  assign _GEN_6399 = {{16'd0}, _T_24414};
  assign _T_53519 = _GEN_6399 << 16;
  assign _GEN_6400 = {{8'd0}, _T_53483};
  assign _T_53523 = _GEN_6400 | _T_53519;
  assign _GEN_6401 = {{24'd0}, _T_24416};
  assign _T_53559 = _GEN_6401 << 24;
  assign _GEN_6402 = {{8'd0}, _T_53523};
  assign _T_53563 = _GEN_6402 | _T_53559;
  assign _GEN_6403 = {{8'd0}, _T_25508};
  assign _T_53639 = _GEN_6403 << 8;
  assign _GEN_6404 = {{8'd0}, _T_25506};
  assign _T_53643 = _GEN_6404 | _T_53639;
  assign _GEN_6405 = {{16'd0}, _T_25510};
  assign _T_53679 = _GEN_6405 << 16;
  assign _GEN_6406 = {{8'd0}, _T_53643};
  assign _T_53683 = _GEN_6406 | _T_53679;
  assign _GEN_6407 = {{24'd0}, _T_25512};
  assign _T_53719 = _GEN_6407 << 24;
  assign _GEN_6408 = {{8'd0}, _T_53683};
  assign _T_53723 = _GEN_6408 | _T_53719;
  assign _GEN_6409 = {{8'd0}, _T_25612};
  assign _T_53959 = _GEN_6409 << 8;
  assign _GEN_6410 = {{8'd0}, _T_25610};
  assign _T_53963 = _GEN_6410 | _T_53959;
  assign _GEN_6411 = {{16'd0}, _T_25614};
  assign _T_53999 = _GEN_6411 << 16;
  assign _GEN_6412 = {{8'd0}, _T_53963};
  assign _T_54003 = _GEN_6412 | _T_53999;
  assign _GEN_6413 = {{24'd0}, _T_25616};
  assign _T_54039 = _GEN_6413 << 24;
  assign _GEN_6414 = {{8'd0}, _T_54003};
  assign _T_54043 = _GEN_6414 | _T_54039;
  assign _T_54063 = _T_99458 & _T_35050;
  assign _GEN_2464 = _T_54063 ? _T_35064 : _GEN_337;
  assign _T_54103 = _T_99458 & _T_35090;
  assign _GEN_2465 = _T_54103 ? _T_35104 : _GEN_338;
  assign _T_54143 = _T_99458 & _T_35130;
  assign _GEN_2466 = _T_54143 ? _T_35144 : _GEN_339;
  assign _T_54183 = _T_99458 & _T_35170;
  assign _GEN_2467 = _T_54183 ? _T_35184 : _GEN_340;
  assign _GEN_6421 = {{8'd0}, _T_24844};
  assign _T_54279 = _GEN_6421 << 8;
  assign _GEN_6422 = {{8'd0}, _T_24842};
  assign _T_54283 = _GEN_6422 | _T_54279;
  assign _GEN_6423 = {{16'd0}, _T_24846};
  assign _T_54319 = _GEN_6423 << 16;
  assign _GEN_6424 = {{8'd0}, _T_54283};
  assign _T_54323 = _GEN_6424 | _T_54319;
  assign _GEN_6425 = {{24'd0}, _T_24848};
  assign _T_54359 = _GEN_6425 << 24;
  assign _GEN_6426 = {{8'd0}, _T_54323};
  assign _T_54363 = _GEN_6426 | _T_54359;
  assign _GEN_6427 = {{8'd0}, _T_25356};
  assign _T_54599 = _GEN_6427 << 8;
  assign _GEN_6428 = {{8'd0}, _T_25354};
  assign _T_54603 = _GEN_6428 | _T_54599;
  assign _GEN_6429 = {{16'd0}, _T_25358};
  assign _T_54639 = _GEN_6429 << 16;
  assign _GEN_6430 = {{8'd0}, _T_54603};
  assign _T_54643 = _GEN_6430 | _T_54639;
  assign _GEN_6431 = {{24'd0}, _T_25360};
  assign _T_54679 = _GEN_6431 << 24;
  assign _GEN_6432 = {{8'd0}, _T_54643};
  assign _T_54683 = _GEN_6432 | _T_54679;
  assign _GEN_6433 = {{8'd0}, _T_24668};
  assign _T_54759 = _GEN_6433 << 8;
  assign _GEN_6434 = {{8'd0}, _T_24666};
  assign _T_54763 = _GEN_6434 | _T_54759;
  assign _GEN_6435 = {{16'd0}, _T_24670};
  assign _T_54799 = _GEN_6435 << 16;
  assign _GEN_6436 = {{8'd0}, _T_54763};
  assign _T_54803 = _GEN_6436 | _T_54799;
  assign _GEN_6437 = {{24'd0}, _T_24672};
  assign _T_54839 = _GEN_6437 << 24;
  assign _GEN_6438 = {{8'd0}, _T_54803};
  assign _T_54843 = _GEN_6438 | _T_54839;
  assign _GEN_6439 = {{8'd0}, _T_25724};
  assign _T_54919 = _GEN_6439 << 8;
  assign _GEN_6440 = {{8'd0}, _T_25722};
  assign _T_54923 = _GEN_6440 | _T_54919;
  assign _GEN_6441 = {{16'd0}, _T_25726};
  assign _T_54959 = _GEN_6441 << 16;
  assign _GEN_6442 = {{8'd0}, _T_54923};
  assign _T_54963 = _GEN_6442 | _T_54959;
  assign _GEN_6443 = {{24'd0}, _T_25728};
  assign _T_54999 = _GEN_6443 << 24;
  assign _GEN_6444 = {{8'd0}, _T_54963};
  assign _T_55003 = _GEN_6444 | _T_54999;
  assign _GEN_6445 = {{8'd0}, _T_24444};
  assign _T_55079 = _GEN_6445 << 8;
  assign _GEN_6446 = {{8'd0}, _T_24442};
  assign _T_55083 = _GEN_6446 | _T_55079;
  assign _GEN_6447 = {{16'd0}, _T_24446};
  assign _T_55119 = _GEN_6447 << 16;
  assign _GEN_6448 = {{8'd0}, _T_55083};
  assign _T_55123 = _GEN_6448 | _T_55119;
  assign _GEN_6449 = {{24'd0}, _T_24448};
  assign _T_55159 = _GEN_6449 << 24;
  assign _GEN_6450 = {{8'd0}, _T_55123};
  assign _T_55163 = _GEN_6450 | _T_55159;
  assign _GEN_6451 = {{8'd0}, _T_23828};
  assign _T_55239 = _GEN_6451 << 8;
  assign _GEN_6452 = {{8'd0}, _T_23826};
  assign _T_55243 = _GEN_6452 | _T_55239;
  assign _GEN_6453 = {{16'd0}, _T_23830};
  assign _T_55279 = _GEN_6453 << 16;
  assign _GEN_6454 = {{8'd0}, _T_55243};
  assign _T_55283 = _GEN_6454 | _T_55279;
  assign _GEN_6455 = {{24'd0}, _T_23832};
  assign _T_55319 = _GEN_6455 << 24;
  assign _GEN_6456 = {{8'd0}, _T_55283};
  assign _T_55323 = _GEN_6456 | _T_55319;
  assign _GEN_6457 = {{8'd0}, _T_24580};
  assign _T_55399 = _GEN_6457 << 8;
  assign _GEN_6458 = {{8'd0}, _T_24578};
  assign _T_55403 = _GEN_6458 | _T_55399;
  assign _GEN_6459 = {{16'd0}, _T_24582};
  assign _T_55439 = _GEN_6459 << 16;
  assign _GEN_6460 = {{8'd0}, _T_55403};
  assign _T_55443 = _GEN_6460 | _T_55439;
  assign _GEN_6461 = {{24'd0}, _T_24584};
  assign _T_55479 = _GEN_6461 << 24;
  assign _GEN_6462 = {{8'd0}, _T_55443};
  assign _T_55483 = _GEN_6462 | _T_55479;
  assign _GEN_6463 = {{8'd0}, _T_25764};
  assign _T_55559 = _GEN_6463 << 8;
  assign _GEN_6464 = {{8'd0}, _T_25762};
  assign _T_55563 = _GEN_6464 | _T_55559;
  assign _GEN_6465 = {{16'd0}, _T_25766};
  assign _T_55599 = _GEN_6465 << 16;
  assign _GEN_6466 = {{8'd0}, _T_55563};
  assign _T_55603 = _GEN_6466 | _T_55599;
  assign _GEN_6467 = {{24'd0}, _T_25768};
  assign _T_55639 = _GEN_6467 << 24;
  assign _GEN_6468 = {{8'd0}, _T_55603};
  assign _T_55643 = _GEN_6468 | _T_55639;
  assign _GEN_6469 = {{8'd0}, _T_24188};
  assign _T_55719 = _GEN_6469 << 8;
  assign _GEN_6470 = {{8'd0}, _T_24186};
  assign _T_55723 = _GEN_6470 | _T_55719;
  assign _GEN_6471 = {{16'd0}, _T_24190};
  assign _T_55759 = _GEN_6471 << 16;
  assign _GEN_6472 = {{8'd0}, _T_55723};
  assign _T_55763 = _GEN_6472 | _T_55759;
  assign _GEN_6473 = {{24'd0}, _T_24192};
  assign _T_55799 = _GEN_6473 << 24;
  assign _GEN_6474 = {{8'd0}, _T_55763};
  assign _T_55803 = _GEN_6474 | _T_55799;
  assign _GEN_6475 = {{8'd0}, _T_24884};
  assign _T_55879 = _GEN_6475 << 8;
  assign _GEN_6476 = {{8'd0}, _T_24882};
  assign _T_55883 = _GEN_6476 | _T_55879;
  assign _GEN_6477 = {{16'd0}, _T_24886};
  assign _T_55919 = _GEN_6477 << 16;
  assign _GEN_6478 = {{8'd0}, _T_55883};
  assign _T_55923 = _GEN_6478 | _T_55919;
  assign _GEN_6479 = {{24'd0}, _T_24888};
  assign _T_55959 = _GEN_6479 << 24;
  assign _GEN_6480 = {{8'd0}, _T_55923};
  assign _T_55963 = _GEN_6480 | _T_55959;
  assign _GEN_6481 = {{8'd0}, _T_24084};
  assign _T_56199 = _GEN_6481 << 8;
  assign _GEN_6482 = {{8'd0}, _T_24082};
  assign _T_56203 = _GEN_6482 | _T_56199;
  assign _GEN_6483 = {{16'd0}, _T_24086};
  assign _T_56239 = _GEN_6483 << 16;
  assign _GEN_6484 = {{8'd0}, _T_56203};
  assign _T_56243 = _GEN_6484 | _T_56239;
  assign _GEN_6485 = {{24'd0}, _T_24088};
  assign _T_56279 = _GEN_6485 << 24;
  assign _GEN_6486 = {{8'd0}, _T_56243};
  assign _T_56283 = _GEN_6486 | _T_56279;
  assign _GEN_6487 = {{8'd0}, _T_24996};
  assign _T_56359 = _GEN_6487 << 8;
  assign _GEN_6488 = {{8'd0}, _T_24994};
  assign _T_56363 = _GEN_6488 | _T_56359;
  assign _GEN_6489 = {{16'd0}, _T_24998};
  assign _T_56399 = _GEN_6489 << 16;
  assign _GEN_6490 = {{8'd0}, _T_56363};
  assign _T_56403 = _GEN_6490 | _T_56399;
  assign _GEN_6491 = {{24'd0}, _T_25000};
  assign _T_56439 = _GEN_6491 << 24;
  assign _GEN_6492 = {{8'd0}, _T_56403};
  assign _T_56443 = _GEN_6492 | _T_56439;
  assign _GEN_6493 = {{8'd0}, _T_25100};
  assign _T_56519 = _GEN_6493 << 8;
  assign _GEN_6494 = {{8'd0}, _T_25098};
  assign _T_56523 = _GEN_6494 | _T_56519;
  assign _GEN_6495 = {{16'd0}, _T_25102};
  assign _T_56559 = _GEN_6495 << 16;
  assign _GEN_6496 = {{8'd0}, _T_56523};
  assign _T_56563 = _GEN_6496 | _T_56559;
  assign _GEN_6497 = {{24'd0}, _T_25104};
  assign _T_56599 = _GEN_6497 << 24;
  assign _GEN_6498 = {{8'd0}, _T_56563};
  assign _T_56603 = _GEN_6498 | _T_56599;
  assign _GEN_6499 = {{8'd0}, _T_25140};
  assign _T_56839 = _GEN_6499 << 8;
  assign _GEN_6500 = {{8'd0}, _T_25138};
  assign _T_56843 = _GEN_6500 | _T_56839;
  assign _GEN_6501 = {{16'd0}, _T_25142};
  assign _T_56879 = _GEN_6501 << 16;
  assign _GEN_6502 = {{8'd0}, _T_56843};
  assign _T_56883 = _GEN_6502 | _T_56879;
  assign _GEN_6503 = {{24'd0}, _T_25144};
  assign _T_56919 = _GEN_6503 << 24;
  assign _GEN_6504 = {{8'd0}, _T_56883};
  assign _T_56923 = _GEN_6504 | _T_56919;
  assign _GEN_6505 = {{8'd0}, _T_23812};
  assign _T_56999 = _GEN_6505 << 8;
  assign _GEN_6506 = {{8'd0}, _T_23810};
  assign _T_57003 = _GEN_6506 | _T_56999;
  assign _GEN_6507 = {{16'd0}, _T_23814};
  assign _T_57039 = _GEN_6507 << 16;
  assign _GEN_6508 = {{8'd0}, _T_57003};
  assign _T_57043 = _GEN_6508 | _T_57039;
  assign _GEN_6509 = {{24'd0}, _T_23816};
  assign _T_57079 = _GEN_6509 << 24;
  assign _GEN_6510 = {{8'd0}, _T_57043};
  assign _T_57083 = _GEN_6510 | _T_57079;
  assign _GEN_6511 = {{8'd0}, _T_23932};
  assign _T_57159 = _GEN_6511 << 8;
  assign _GEN_6512 = {{8'd0}, _T_23930};
  assign _T_57163 = _GEN_6512 | _T_57159;
  assign _GEN_6513 = {{16'd0}, _T_23934};
  assign _T_57199 = _GEN_6513 << 16;
  assign _GEN_6514 = {{8'd0}, _T_57163};
  assign _T_57203 = _GEN_6514 | _T_57199;
  assign _GEN_6515 = {{24'd0}, _T_23936};
  assign _T_57239 = _GEN_6515 << 24;
  assign _GEN_6516 = {{8'd0}, _T_57203};
  assign _T_57243 = _GEN_6516 | _T_57239;
  assign _T_57263 = _T_98274 & _T_50170;
  assign _T_57264 = io_hart_in_0_a_bits_data[9:0];
  assign _GEN_6517 = {{8'd0}, _T_24068};
  assign _T_57359 = _GEN_6517 << 8;
  assign _GEN_6518 = {{8'd0}, _T_24066};
  assign _T_57363 = _GEN_6518 | _T_57359;
  assign _GEN_6519 = {{16'd0}, _T_24070};
  assign _T_57399 = _GEN_6519 << 16;
  assign _GEN_6520 = {{8'd0}, _T_57363};
  assign _T_57403 = _GEN_6520 | _T_57399;
  assign _GEN_6521 = {{24'd0}, _T_24072};
  assign _T_57439 = _GEN_6521 << 24;
  assign _GEN_6522 = {{8'd0}, _T_57403};
  assign _T_57443 = _GEN_6522 | _T_57439;
  assign _GEN_6523 = {{8'd0}, _T_25252};
  assign _T_57519 = _GEN_6523 << 8;
  assign _GEN_6524 = {{8'd0}, _T_25250};
  assign _T_57523 = _GEN_6524 | _T_57519;
  assign _GEN_6525 = {{16'd0}, _T_25254};
  assign _T_57559 = _GEN_6525 << 16;
  assign _GEN_6526 = {{8'd0}, _T_57523};
  assign _T_57563 = _GEN_6526 | _T_57559;
  assign _GEN_6527 = {{24'd0}, _T_25256};
  assign _T_57599 = _GEN_6527 << 24;
  assign _GEN_6528 = {{8'd0}, _T_57563};
  assign _T_57603 = _GEN_6528 | _T_57599;
  assign _GEN_6529 = {{8'd0}, _T_24700};
  assign _T_57679 = _GEN_6529 << 8;
  assign _GEN_6530 = {{8'd0}, _T_24698};
  assign _T_57683 = _GEN_6530 | _T_57679;
  assign _GEN_6531 = {{16'd0}, _T_24702};
  assign _T_57719 = _GEN_6531 << 16;
  assign _GEN_6532 = {{8'd0}, _T_57683};
  assign _T_57723 = _GEN_6532 | _T_57719;
  assign _GEN_6533 = {{24'd0}, _T_24704};
  assign _T_57759 = _GEN_6533 << 24;
  assign _GEN_6534 = {{8'd0}, _T_57723};
  assign _T_57763 = _GEN_6534 | _T_57759;
  assign _GEN_6535 = {{8'd0}, _T_25084};
  assign _T_57839 = _GEN_6535 << 8;
  assign _GEN_6536 = {{8'd0}, _T_25082};
  assign _T_57843 = _GEN_6536 | _T_57839;
  assign _GEN_6537 = {{16'd0}, _T_25086};
  assign _T_57879 = _GEN_6537 << 16;
  assign _GEN_6538 = {{8'd0}, _T_57843};
  assign _T_57883 = _GEN_6538 | _T_57879;
  assign _GEN_6539 = {{24'd0}, _T_25088};
  assign _T_57919 = _GEN_6539 << 24;
  assign _GEN_6540 = {{8'd0}, _T_57883};
  assign _T_57923 = _GEN_6540 | _T_57919;
  assign _GEN_6541 = {{8'd0}, _T_24916};
  assign _T_57999 = _GEN_6541 << 8;
  assign _GEN_6542 = {{8'd0}, _T_24914};
  assign _T_58003 = _GEN_6542 | _T_57999;
  assign _GEN_6543 = {{16'd0}, _T_24918};
  assign _T_58039 = _GEN_6543 << 16;
  assign _GEN_6544 = {{8'd0}, _T_58003};
  assign _T_58043 = _GEN_6544 | _T_58039;
  assign _GEN_6545 = {{24'd0}, _T_24920};
  assign _T_58079 = _GEN_6545 << 24;
  assign _GEN_6546 = {{8'd0}, _T_58043};
  assign _T_58083 = _GEN_6546 | _T_58079;
  assign _GEN_6547 = {{8'd0}, _T_23988};
  assign _T_58159 = _GEN_6547 << 8;
  assign _GEN_6548 = {{8'd0}, _T_23986};
  assign _T_58163 = _GEN_6548 | _T_58159;
  assign _GEN_6549 = {{16'd0}, _T_23990};
  assign _T_58199 = _GEN_6549 << 16;
  assign _GEN_6550 = {{8'd0}, _T_58163};
  assign _T_58203 = _GEN_6550 | _T_58199;
  assign _GEN_6551 = {{24'd0}, _T_23992};
  assign _T_58239 = _GEN_6551 << 24;
  assign _GEN_6552 = {{8'd0}, _T_58203};
  assign _T_58243 = _GEN_6552 | _T_58239;
  assign _GEN_6553 = {{8'd0}, _T_24028};
  assign _T_58319 = _GEN_6553 << 8;
  assign _GEN_6554 = {{8'd0}, _T_24026};
  assign _T_58323 = _GEN_6554 | _T_58319;
  assign _GEN_6555 = {{16'd0}, _T_24030};
  assign _T_58359 = _GEN_6555 << 16;
  assign _GEN_6556 = {{8'd0}, _T_58323};
  assign _T_58363 = _GEN_6556 | _T_58359;
  assign _GEN_6557 = {{24'd0}, _T_24032};
  assign _T_58399 = _GEN_6557 << 24;
  assign _GEN_6558 = {{8'd0}, _T_58363};
  assign _T_58403 = _GEN_6558 | _T_58399;
  assign _GEN_6559 = {{8'd0}, _T_23948};
  assign _T_58479 = _GEN_6559 << 8;
  assign _GEN_6560 = {{8'd0}, _T_23946};
  assign _T_58483 = _GEN_6560 | _T_58479;
  assign _GEN_6561 = {{16'd0}, _T_23950};
  assign _T_58519 = _GEN_6561 << 16;
  assign _GEN_6562 = {{8'd0}, _T_58483};
  assign _T_58523 = _GEN_6562 | _T_58519;
  assign _GEN_6563 = {{24'd0}, _T_23952};
  assign _T_58559 = _GEN_6563 << 24;
  assign _GEN_6564 = {{8'd0}, _T_58523};
  assign _T_58563 = _GEN_6564 | _T_58559;
  assign _GEN_6565 = {{8'd0}, _T_23772};
  assign _T_58639 = _GEN_6565 << 8;
  assign _GEN_6566 = {{8'd0}, _T_23770};
  assign _T_58643 = _GEN_6566 | _T_58639;
  assign _GEN_6567 = {{16'd0}, _T_23774};
  assign _T_58679 = _GEN_6567 << 16;
  assign _GEN_6568 = {{8'd0}, _T_58643};
  assign _T_58683 = _GEN_6568 | _T_58679;
  assign _GEN_6569 = {{24'd0}, _T_23776};
  assign _T_58719 = _GEN_6569 << 24;
  assign _GEN_6570 = {{8'd0}, _T_58683};
  assign _T_58723 = _GEN_6570 | _T_58719;
  assign _GEN_6571 = {{8'd0}, _T_25004};
  assign _T_58799 = _GEN_6571 << 8;
  assign _GEN_6572 = {{8'd0}, _T_25002};
  assign _T_58803 = _GEN_6572 | _T_58799;
  assign _GEN_6573 = {{16'd0}, _T_25006};
  assign _T_58839 = _GEN_6573 << 16;
  assign _GEN_6574 = {{8'd0}, _T_58803};
  assign _T_58843 = _GEN_6574 | _T_58839;
  assign _GEN_6575 = {{24'd0}, _T_25008};
  assign _T_58879 = _GEN_6575 << 24;
  assign _GEN_6576 = {{8'd0}, _T_58843};
  assign _T_58883 = _GEN_6576 | _T_58879;
  assign _GEN_6577 = {{8'd0}, _T_24828};
  assign _T_58959 = _GEN_6577 << 8;
  assign _GEN_6578 = {{8'd0}, _T_24826};
  assign _T_58963 = _GEN_6578 | _T_58959;
  assign _GEN_6579 = {{16'd0}, _T_24830};
  assign _T_58999 = _GEN_6579 << 16;
  assign _GEN_6580 = {{8'd0}, _T_58963};
  assign _T_59003 = _GEN_6580 | _T_58999;
  assign _GEN_6581 = {{24'd0}, _T_24832};
  assign _T_59039 = _GEN_6581 << 24;
  assign _GEN_6582 = {{8'd0}, _T_59003};
  assign _T_59043 = _GEN_6582 | _T_59039;
  assign _GEN_6583 = {{8'd0}, _T_25260};
  assign _T_59119 = _GEN_6583 << 8;
  assign _GEN_6584 = {{8'd0}, _T_25258};
  assign _T_59123 = _GEN_6584 | _T_59119;
  assign _GEN_6585 = {{16'd0}, _T_25262};
  assign _T_59159 = _GEN_6585 << 16;
  assign _GEN_6586 = {{8'd0}, _T_59123};
  assign _T_59163 = _GEN_6586 | _T_59159;
  assign _GEN_6587 = {{24'd0}, _T_25264};
  assign _T_59199 = _GEN_6587 << 24;
  assign _GEN_6588 = {{8'd0}, _T_59163};
  assign _T_59203 = _GEN_6588 | _T_59199;
  assign _GEN_6589 = {{8'd0}, _T_24756};
  assign _T_59279 = _GEN_6589 << 8;
  assign _GEN_6590 = {{8'd0}, _T_24754};
  assign _T_59283 = _GEN_6590 | _T_59279;
  assign _GEN_6591 = {{16'd0}, _T_24758};
  assign _T_59319 = _GEN_6591 << 16;
  assign _GEN_6592 = {{8'd0}, _T_59283};
  assign _T_59323 = _GEN_6592 | _T_59319;
  assign _GEN_6593 = {{24'd0}, _T_24760};
  assign _T_59359 = _GEN_6593 << 24;
  assign _GEN_6594 = {{8'd0}, _T_59323};
  assign _T_59363 = _GEN_6594 | _T_59359;
  assign _GEN_6595 = {{8'd0}, _T_24204};
  assign _T_59439 = _GEN_6595 << 8;
  assign _GEN_6596 = {{8'd0}, _T_24202};
  assign _T_59443 = _GEN_6596 | _T_59439;
  assign _GEN_6597 = {{16'd0}, _T_24206};
  assign _T_59479 = _GEN_6597 << 16;
  assign _GEN_6598 = {{8'd0}, _T_59443};
  assign _T_59483 = _GEN_6598 | _T_59479;
  assign _GEN_6599 = {{24'd0}, _T_24208};
  assign _T_59519 = _GEN_6599 << 24;
  assign _GEN_6600 = {{8'd0}, _T_59483};
  assign _T_59523 = _GEN_6600 | _T_59519;
  assign _GEN_6601 = {{8'd0}, _T_25684};
  assign _T_59599 = _GEN_6601 << 8;
  assign _GEN_6602 = {{8'd0}, _T_25682};
  assign _T_59603 = _GEN_6602 | _T_59599;
  assign _GEN_6603 = {{16'd0}, _T_25686};
  assign _T_59639 = _GEN_6603 << 16;
  assign _GEN_6604 = {{8'd0}, _T_59603};
  assign _T_59643 = _GEN_6604 | _T_59639;
  assign _GEN_6605 = {{24'd0}, _T_25688};
  assign _T_59679 = _GEN_6605 << 24;
  assign _GEN_6606 = {{8'd0}, _T_59643};
  assign _T_59683 = _GEN_6606 | _T_59679;
  assign _GEN_6607 = {{8'd0}, _T_25428};
  assign _T_59759 = _GEN_6607 << 8;
  assign _GEN_6608 = {{8'd0}, _T_25426};
  assign _T_59763 = _GEN_6608 | _T_59759;
  assign _GEN_6609 = {{16'd0}, _T_25430};
  assign _T_59799 = _GEN_6609 << 16;
  assign _GEN_6610 = {{8'd0}, _T_59763};
  assign _T_59803 = _GEN_6610 | _T_59799;
  assign _GEN_6611 = {{24'd0}, _T_25432};
  assign _T_59839 = _GEN_6611 << 24;
  assign _GEN_6612 = {{8'd0}, _T_59803};
  assign _T_59843 = _GEN_6612 | _T_59839;
  assign _GEN_6613 = {{8'd0}, _T_24380};
  assign _T_59919 = _GEN_6613 << 8;
  assign _GEN_6614 = {{8'd0}, _T_24378};
  assign _T_59923 = _GEN_6614 | _T_59919;
  assign _GEN_6615 = {{16'd0}, _T_24382};
  assign _T_59959 = _GEN_6615 << 16;
  assign _GEN_6616 = {{8'd0}, _T_59923};
  assign _T_59963 = _GEN_6616 | _T_59959;
  assign _GEN_6617 = {{24'd0}, _T_24384};
  assign _T_59999 = _GEN_6617 << 24;
  assign _GEN_6618 = {{8'd0}, _T_59963};
  assign _T_60003 = _GEN_6618 | _T_59999;
  assign _GEN_6619 = {{8'd0}, _T_24500};
  assign _T_60079 = _GEN_6619 << 8;
  assign _GEN_6620 = {{8'd0}, _T_24498};
  assign _T_60083 = _GEN_6620 | _T_60079;
  assign _GEN_6621 = {{16'd0}, _T_24502};
  assign _T_60119 = _GEN_6621 << 16;
  assign _GEN_6622 = {{8'd0}, _T_60083};
  assign _T_60123 = _GEN_6622 | _T_60119;
  assign _GEN_6623 = {{24'd0}, _T_24504};
  assign _T_60159 = _GEN_6623 << 24;
  assign _GEN_6624 = {{8'd0}, _T_60123};
  assign _T_60163 = _GEN_6624 | _T_60159;
  assign _GEN_6625 = {{8'd0}, _T_24948};
  assign _T_60239 = _GEN_6625 << 8;
  assign _GEN_6626 = {{8'd0}, _T_24946};
  assign _T_60243 = _GEN_6626 | _T_60239;
  assign _GEN_6627 = {{16'd0}, _T_24950};
  assign _T_60279 = _GEN_6627 << 16;
  assign _GEN_6628 = {{8'd0}, _T_60243};
  assign _T_60283 = _GEN_6628 | _T_60279;
  assign _GEN_6629 = {{24'd0}, _T_24952};
  assign _T_60319 = _GEN_6629 << 24;
  assign _GEN_6630 = {{8'd0}, _T_60283};
  assign _T_60323 = _GEN_6630 | _T_60319;
  assign _T_60343 = _T_99514 & _T_35050;
  assign _GEN_2469 = _T_60343 ? _T_35064 : _GEN_365;
  assign _T_60383 = _T_99514 & _T_35090;
  assign _GEN_2470 = _T_60383 ? _T_35104 : _GEN_366;
  assign _T_60423 = _T_99514 & _T_35130;
  assign _GEN_2471 = _T_60423 ? _T_35144 : _GEN_367;
  assign _T_60463 = _T_99514 & _T_35170;
  assign _GEN_2472 = _T_60463 ? _T_35184 : _GEN_368;
  assign _GEN_6637 = {{8'd0}, _T_23892};
  assign _T_60559 = _GEN_6637 << 8;
  assign _GEN_6638 = {{8'd0}, _T_23890};
  assign _T_60563 = _GEN_6638 | _T_60559;
  assign _GEN_6639 = {{16'd0}, _T_23894};
  assign _T_60599 = _GEN_6639 << 16;
  assign _GEN_6640 = {{8'd0}, _T_60563};
  assign _T_60603 = _GEN_6640 | _T_60599;
  assign _GEN_6641 = {{24'd0}, _T_23896};
  assign _T_60639 = _GEN_6641 << 24;
  assign _GEN_6642 = {{8'd0}, _T_60603};
  assign _T_60643 = _GEN_6642 | _T_60639;
  assign _GEN_6643 = {{8'd0}, _T_25052};
  assign _T_60719 = _GEN_6643 << 8;
  assign _GEN_6644 = {{8'd0}, _T_25050};
  assign _T_60723 = _GEN_6644 | _T_60719;
  assign _GEN_6645 = {{16'd0}, _T_25054};
  assign _T_60759 = _GEN_6645 << 16;
  assign _GEN_6646 = {{8'd0}, _T_60723};
  assign _T_60763 = _GEN_6646 | _T_60759;
  assign _GEN_6647 = {{24'd0}, _T_25056};
  assign _T_60799 = _GEN_6647 << 24;
  assign _GEN_6648 = {{8'd0}, _T_60763};
  assign _T_60803 = _GEN_6648 | _T_60799;
  assign _GEN_6649 = {{8'd0}, _T_24716};
  assign _T_60879 = _GEN_6649 << 8;
  assign _GEN_6650 = {{8'd0}, _T_24714};
  assign _T_60883 = _GEN_6650 | _T_60879;
  assign _GEN_6651 = {{16'd0}, _T_24718};
  assign _T_60919 = _GEN_6651 << 16;
  assign _GEN_6652 = {{8'd0}, _T_60883};
  assign _T_60923 = _GEN_6652 | _T_60919;
  assign _GEN_6653 = {{24'd0}, _T_24720};
  assign _T_60959 = _GEN_6653 << 24;
  assign _GEN_6654 = {{8'd0}, _T_60923};
  assign _T_60963 = _GEN_6654 | _T_60959;
  assign _GEN_6655 = {{8'd0}, _T_24596};
  assign _T_61039 = _GEN_6655 << 8;
  assign _GEN_6656 = {{8'd0}, _T_24594};
  assign _T_61043 = _GEN_6656 | _T_61039;
  assign _GEN_6657 = {{16'd0}, _T_24598};
  assign _T_61079 = _GEN_6657 << 16;
  assign _GEN_6658 = {{8'd0}, _T_61043};
  assign _T_61083 = _GEN_6658 | _T_61079;
  assign _GEN_6659 = {{24'd0}, _T_24600};
  assign _T_61119 = _GEN_6659 << 24;
  assign _GEN_6660 = {{8'd0}, _T_61083};
  assign _T_61123 = _GEN_6660 | _T_61119;
  assign _GEN_6661 = {{8'd0}, _T_25308};
  assign _T_61199 = _GEN_6661 << 8;
  assign _GEN_6662 = {{8'd0}, _T_25306};
  assign _T_61203 = _GEN_6662 | _T_61199;
  assign _GEN_6663 = {{16'd0}, _T_25310};
  assign _T_61239 = _GEN_6663 << 16;
  assign _GEN_6664 = {{8'd0}, _T_61203};
  assign _T_61243 = _GEN_6664 | _T_61239;
  assign _GEN_6665 = {{24'd0}, _T_25312};
  assign _T_61279 = _GEN_6665 << 24;
  assign _GEN_6666 = {{8'd0}, _T_61243};
  assign _T_61283 = _GEN_6666 | _T_61279;
  assign _GEN_6667 = {{8'd0}, _T_24244};
  assign _T_61359 = _GEN_6667 << 8;
  assign _GEN_6668 = {{8'd0}, _T_24242};
  assign _T_61363 = _GEN_6668 | _T_61359;
  assign _GEN_6669 = {{16'd0}, _T_24246};
  assign _T_61399 = _GEN_6669 << 16;
  assign _GEN_6670 = {{8'd0}, _T_61363};
  assign _T_61403 = _GEN_6670 | _T_61399;
  assign _GEN_6671 = {{24'd0}, _T_24248};
  assign _T_61439 = _GEN_6671 << 24;
  assign _GEN_6672 = {{8'd0}, _T_61403};
  assign _T_61443 = _GEN_6672 | _T_61439;
  assign _GEN_6673 = {{8'd0}, _T_25772};
  assign _T_61519 = _GEN_6673 << 8;
  assign _GEN_6674 = {{8'd0}, _T_25770};
  assign _T_61523 = _GEN_6674 | _T_61519;
  assign _GEN_6675 = {{16'd0}, _T_25774};
  assign _T_61559 = _GEN_6675 << 16;
  assign _GEN_6676 = {{8'd0}, _T_61523};
  assign _T_61563 = _GEN_6676 | _T_61559;
  assign _GEN_6677 = {{24'd0}, _T_25776};
  assign _T_61599 = _GEN_6677 << 24;
  assign _GEN_6678 = {{8'd0}, _T_61563};
  assign _T_61603 = _GEN_6678 | _T_61599;
  assign _GEN_6679 = {{8'd0}, _T_25172};
  assign _T_61679 = _GEN_6679 << 8;
  assign _GEN_6680 = {{8'd0}, _T_25170};
  assign _T_61683 = _GEN_6680 | _T_61679;
  assign _GEN_6681 = {{16'd0}, _T_25174};
  assign _T_61719 = _GEN_6681 << 16;
  assign _GEN_6682 = {{8'd0}, _T_61683};
  assign _T_61723 = _GEN_6682 | _T_61719;
  assign _GEN_6683 = {{24'd0}, _T_25176};
  assign _T_61759 = _GEN_6683 << 24;
  assign _GEN_6684 = {{8'd0}, _T_61723};
  assign _T_61763 = _GEN_6684 | _T_61759;
  assign _GEN_6685 = {{8'd0}, _T_24124};
  assign _T_61839 = _GEN_6685 << 8;
  assign _GEN_6686 = {{8'd0}, _T_24122};
  assign _T_61843 = _GEN_6686 | _T_61839;
  assign _GEN_6687 = {{16'd0}, _T_24126};
  assign _T_61879 = _GEN_6687 << 16;
  assign _GEN_6688 = {{8'd0}, _T_61843};
  assign _T_61883 = _GEN_6688 | _T_61879;
  assign _GEN_6689 = {{24'd0}, _T_24128};
  assign _T_61919 = _GEN_6689 << 24;
  assign _GEN_6690 = {{8'd0}, _T_61883};
  assign _T_61923 = _GEN_6690 | _T_61919;
  assign _GEN_6691 = {{8'd0}, _T_23868};
  assign _T_61999 = _GEN_6691 << 8;
  assign _GEN_6692 = {{8'd0}, _T_23866};
  assign _T_62003 = _GEN_6692 | _T_61999;
  assign _GEN_6693 = {{16'd0}, _T_23870};
  assign _T_62039 = _GEN_6693 << 16;
  assign _GEN_6694 = {{8'd0}, _T_62003};
  assign _T_62043 = _GEN_6694 | _T_62039;
  assign _GEN_6695 = {{24'd0}, _T_23872};
  assign _T_62079 = _GEN_6695 << 24;
  assign _GEN_6696 = {{8'd0}, _T_62043};
  assign _T_62083 = _GEN_6696 | _T_62079;
  assign _T_62103 = _T_99426 & _T_35050;
  assign _GEN_2473 = _T_62103 ? _T_35064 : _GEN_321;
  assign _T_62143 = _T_99426 & _T_35090;
  assign _GEN_2474 = _T_62143 ? _T_35104 : _GEN_322;
  assign _T_62183 = _T_99426 & _T_35130;
  assign _GEN_2475 = _T_62183 ? _T_35144 : _GEN_323;
  assign _T_62223 = _T_99426 & _T_35170;
  assign _GEN_2476 = _T_62223 ? _T_35184 : _GEN_324;
  assign _GEN_6703 = {{8'd0}, _T_25516};
  assign _T_62319 = _GEN_6703 << 8;
  assign _GEN_6704 = {{8'd0}, _T_25514};
  assign _T_62323 = _GEN_6704 | _T_62319;
  assign _GEN_6705 = {{16'd0}, _T_25518};
  assign _T_62359 = _GEN_6705 << 16;
  assign _GEN_6706 = {{8'd0}, _T_62323};
  assign _T_62363 = _GEN_6706 | _T_62359;
  assign _GEN_6707 = {{24'd0}, _T_25520};
  assign _T_62399 = _GEN_6707 << 24;
  assign _GEN_6708 = {{8'd0}, _T_62363};
  assign _T_62403 = _GEN_6708 | _T_62399;
  assign _GEN_6709 = {{8'd0}, _T_24796};
  assign _T_62479 = _GEN_6709 << 8;
  assign _GEN_6710 = {{8'd0}, _T_24794};
  assign _T_62483 = _GEN_6710 | _T_62479;
  assign _GEN_6711 = {{16'd0}, _T_24798};
  assign _T_62519 = _GEN_6711 << 16;
  assign _GEN_6712 = {{8'd0}, _T_62483};
  assign _T_62523 = _GEN_6712 | _T_62519;
  assign _GEN_6713 = {{24'd0}, _T_24800};
  assign _T_62559 = _GEN_6713 << 24;
  assign _GEN_6714 = {{8'd0}, _T_62523};
  assign _T_62563 = _GEN_6714 | _T_62559;
  assign _GEN_6715 = {{8'd0}, _T_25652};
  assign _T_62639 = _GEN_6715 << 8;
  assign _GEN_6716 = {{8'd0}, _T_25650};
  assign _T_62643 = _GEN_6716 | _T_62639;
  assign _GEN_6717 = {{16'd0}, _T_25654};
  assign _T_62679 = _GEN_6717 << 16;
  assign _GEN_6718 = {{8'd0}, _T_62643};
  assign _T_62683 = _GEN_6718 | _T_62679;
  assign _GEN_6719 = {{24'd0}, _T_25656};
  assign _T_62719 = _GEN_6719 << 24;
  assign _GEN_6720 = {{8'd0}, _T_62683};
  assign _T_62723 = _GEN_6720 | _T_62719;
  assign _GEN_6721 = {{8'd0}, _T_24460};
  assign _T_62799 = _GEN_6721 << 8;
  assign _GEN_6722 = {{8'd0}, _T_24458};
  assign _T_62803 = _GEN_6722 | _T_62799;
  assign _GEN_6723 = {{16'd0}, _T_24462};
  assign _T_62839 = _GEN_6723 << 16;
  assign _GEN_6724 = {{8'd0}, _T_62803};
  assign _T_62843 = _GEN_6724 | _T_62839;
  assign _GEN_6725 = {{24'd0}, _T_24464};
  assign _T_62879 = _GEN_6725 << 24;
  assign _GEN_6726 = {{8'd0}, _T_62843};
  assign _T_62883 = _GEN_6726 | _T_62879;
  assign _GEN_6727 = {{8'd0}, _T_24636};
  assign _T_62959 = _GEN_6727 << 8;
  assign _GEN_6728 = {{8'd0}, _T_24634};
  assign _T_62963 = _GEN_6728 | _T_62959;
  assign _GEN_6729 = {{16'd0}, _T_24638};
  assign _T_62999 = _GEN_6729 << 16;
  assign _GEN_6730 = {{8'd0}, _T_62963};
  assign _T_63003 = _GEN_6730 | _T_62999;
  assign _GEN_6731 = {{24'd0}, _T_24640};
  assign _T_63039 = _GEN_6731 << 24;
  assign _GEN_6732 = {{8'd0}, _T_63003};
  assign _T_63043 = _GEN_6732 | _T_63039;
  assign _GEN_6733 = {{8'd0}, _T_24284};
  assign _T_63279 = _GEN_6733 << 8;
  assign _GEN_6734 = {{8'd0}, _T_24282};
  assign _T_63283 = _GEN_6734 | _T_63279;
  assign _GEN_6735 = {{16'd0}, _T_24286};
  assign _T_63319 = _GEN_6735 << 16;
  assign _GEN_6736 = {{8'd0}, _T_63283};
  assign _T_63323 = _GEN_6736 | _T_63319;
  assign _GEN_6737 = {{24'd0}, _T_24288};
  assign _T_63359 = _GEN_6737 << 24;
  assign _GEN_6738 = {{8'd0}, _T_63323};
  assign _T_63363 = _GEN_6738 | _T_63359;
  assign _T_63383 = _T_99466 & _T_35050;
  assign _GEN_2477 = _T_63383 ? _T_35064 : _GEN_341;
  assign _T_63423 = _T_99466 & _T_35090;
  assign _GEN_2478 = _T_63423 ? _T_35104 : _GEN_342;
  assign _T_63463 = _T_99466 & _T_35130;
  assign _GEN_2479 = _T_63463 ? _T_35144 : _GEN_343;
  assign _T_63503 = _T_99466 & _T_35170;
  assign _GEN_2480 = _T_63503 ? _T_35184 : _GEN_344;
  assign _GEN_6745 = {{8'd0}, _T_25564};
  assign _T_63599 = _GEN_6745 << 8;
  assign _GEN_6746 = {{8'd0}, _T_25562};
  assign _T_63603 = _GEN_6746 | _T_63599;
  assign _GEN_6747 = {{16'd0}, _T_25566};
  assign _T_63639 = _GEN_6747 << 16;
  assign _GEN_6748 = {{8'd0}, _T_63603};
  assign _T_63643 = _GEN_6748 | _T_63639;
  assign _GEN_6749 = {{24'd0}, _T_25568};
  assign _T_63679 = _GEN_6749 << 24;
  assign _GEN_6750 = {{8'd0}, _T_63643};
  assign _T_63683 = _GEN_6750 | _T_63679;
  assign _T_63863 = _T_98290 & _T_50170;
  assign _T_63864 = io_hart_in_0_a_bits_data[9:0];
  assign _GEN_6751 = {{8'd0}, _T_24340};
  assign _T_63959 = _GEN_6751 << 8;
  assign _GEN_6752 = {{8'd0}, _T_24338};
  assign _T_63963 = _GEN_6752 | _T_63959;
  assign _GEN_6753 = {{16'd0}, _T_24342};
  assign _T_63999 = _GEN_6753 << 16;
  assign _GEN_6754 = {{8'd0}, _T_63963};
  assign _T_64003 = _GEN_6754 | _T_63999;
  assign _GEN_6755 = {{24'd0}, _T_24344};
  assign _T_64039 = _GEN_6755 << 24;
  assign _GEN_6756 = {{8'd0}, _T_64003};
  assign _T_64043 = _GEN_6756 | _T_64039;
  assign _GEN_6757 = {{8'd0}, _T_25396};
  assign _T_64119 = _GEN_6757 << 8;
  assign _GEN_6758 = {{8'd0}, _T_25394};
  assign _T_64123 = _GEN_6758 | _T_64119;
  assign _GEN_6759 = {{16'd0}, _T_25398};
  assign _T_64159 = _GEN_6759 << 16;
  assign _GEN_6760 = {{8'd0}, _T_64123};
  assign _T_64163 = _GEN_6760 | _T_64159;
  assign _GEN_6761 = {{24'd0}, _T_25400};
  assign _T_64199 = _GEN_6761 << 24;
  assign _GEN_6762 = {{8'd0}, _T_64163};
  assign _T_64203 = _GEN_6762 | _T_64199;
  assign _GEN_6763 = {{8'd0}, _T_24892};
  assign _T_64439 = _GEN_6763 << 8;
  assign _GEN_6764 = {{8'd0}, _T_24890};
  assign _T_64443 = _GEN_6764 | _T_64439;
  assign _GEN_6765 = {{16'd0}, _T_24894};
  assign _T_64479 = _GEN_6765 << 16;
  assign _GEN_6766 = {{8'd0}, _T_64443};
  assign _T_64483 = _GEN_6766 | _T_64479;
  assign _GEN_6767 = {{24'd0}, _T_24896};
  assign _T_64519 = _GEN_6767 << 24;
  assign _GEN_6768 = {{8'd0}, _T_64483};
  assign _T_64523 = _GEN_6768 | _T_64519;
  assign _GEN_6769 = {{8'd0}, _T_23924};
  assign _T_64599 = _GEN_6769 << 8;
  assign _GEN_6770 = {{8'd0}, _T_23922};
  assign _T_64603 = _GEN_6770 | _T_64599;
  assign _GEN_6771 = {{16'd0}, _T_23926};
  assign _T_64639 = _GEN_6771 << 16;
  assign _GEN_6772 = {{8'd0}, _T_64603};
  assign _T_64643 = _GEN_6772 | _T_64639;
  assign _GEN_6773 = {{24'd0}, _T_23928};
  assign _T_64679 = _GEN_6773 << 24;
  assign _GEN_6774 = {{8'd0}, _T_64643};
  assign _T_64683 = _GEN_6774 | _T_64679;
  assign _GEN_6775 = {{8'd0}, _T_25340};
  assign _T_64759 = _GEN_6775 << 8;
  assign _GEN_6776 = {{8'd0}, _T_25338};
  assign _T_64763 = _GEN_6776 | _T_64759;
  assign _GEN_6777 = {{16'd0}, _T_25342};
  assign _T_64799 = _GEN_6777 << 16;
  assign _GEN_6778 = {{8'd0}, _T_64763};
  assign _T_64803 = _GEN_6778 | _T_64799;
  assign _GEN_6779 = {{24'd0}, _T_25344};
  assign _T_64839 = _GEN_6779 << 24;
  assign _GEN_6780 = {{8'd0}, _T_64803};
  assign _T_64843 = _GEN_6780 | _T_64839;
  assign _T_64863 = _T_99546 & _T_35050;
  assign _GEN_2482 = _T_64863 ? _T_35064 : _GEN_381;
  assign _T_64903 = _T_99546 & _T_35090;
  assign _GEN_2483 = _T_64903 ? _T_35104 : _GEN_382;
  assign _T_64943 = _T_99546 & _T_35130;
  assign _GEN_2484 = _T_64943 ? _T_35144 : _GEN_383;
  assign _T_64983 = _T_99546 & _T_35170;
  assign _GEN_2485 = _T_64983 ? _T_35184 : _GEN_384;
  assign _GEN_6787 = {{8'd0}, _T_24852};
  assign _T_65079 = _GEN_6787 << 8;
  assign _GEN_6788 = {{8'd0}, _T_24850};
  assign _T_65083 = _GEN_6788 | _T_65079;
  assign _GEN_6789 = {{16'd0}, _T_24854};
  assign _T_65119 = _GEN_6789 << 16;
  assign _GEN_6790 = {{8'd0}, _T_65083};
  assign _T_65123 = _GEN_6790 | _T_65119;
  assign _GEN_6791 = {{24'd0}, _T_24856};
  assign _T_65159 = _GEN_6791 << 24;
  assign _GEN_6792 = {{8'd0}, _T_65123};
  assign _T_65163 = _GEN_6792 | _T_65159;
  assign _GEN_6793 = {{8'd0}, _T_24148};
  assign _T_65239 = _GEN_6793 << 8;
  assign _GEN_6794 = {{8'd0}, _T_24146};
  assign _T_65243 = _GEN_6794 | _T_65239;
  assign _GEN_6795 = {{16'd0}, _T_24150};
  assign _T_65279 = _GEN_6795 << 16;
  assign _GEN_6796 = {{8'd0}, _T_65243};
  assign _T_65283 = _GEN_6796 | _T_65279;
  assign _GEN_6797 = {{24'd0}, _T_24152};
  assign _T_65319 = _GEN_6797 << 24;
  assign _GEN_6798 = {{8'd0}, _T_65283};
  assign _T_65323 = _GEN_6798 | _T_65319;
  assign _GEN_6799 = {{8'd0}, _T_24092};
  assign _T_65399 = _GEN_6799 << 8;
  assign _GEN_6800 = {{8'd0}, _T_24090};
  assign _T_65403 = _GEN_6800 | _T_65399;
  assign _GEN_6801 = {{16'd0}, _T_24094};
  assign _T_65439 = _GEN_6801 << 16;
  assign _GEN_6802 = {{8'd0}, _T_65403};
  assign _T_65443 = _GEN_6802 | _T_65439;
  assign _GEN_6803 = {{24'd0}, _T_24096};
  assign _T_65479 = _GEN_6803 << 24;
  assign _GEN_6804 = {{8'd0}, _T_65443};
  assign _T_65483 = _GEN_6804 | _T_65479;
  assign _GEN_6805 = {{8'd0}, _T_23836};
  assign _T_65559 = _GEN_6805 << 8;
  assign _GEN_6806 = {{8'd0}, _T_23834};
  assign _T_65563 = _GEN_6806 | _T_65559;
  assign _GEN_6807 = {{16'd0}, _T_23838};
  assign _T_65599 = _GEN_6807 << 16;
  assign _GEN_6808 = {{8'd0}, _T_65563};
  assign _T_65603 = _GEN_6808 | _T_65599;
  assign _GEN_6809 = {{24'd0}, _T_23840};
  assign _T_65639 = _GEN_6809 << 24;
  assign _GEN_6810 = {{8'd0}, _T_65603};
  assign _T_65643 = _GEN_6810 | _T_65639;
  assign _GEN_6811 = {{8'd0}, _T_25740};
  assign _T_65719 = _GEN_6811 << 8;
  assign _GEN_6812 = {{8'd0}, _T_25738};
  assign _T_65723 = _GEN_6812 | _T_65719;
  assign _GEN_6813 = {{16'd0}, _T_25742};
  assign _T_65759 = _GEN_6813 << 16;
  assign _GEN_6814 = {{8'd0}, _T_65723};
  assign _T_65763 = _GEN_6814 | _T_65759;
  assign _GEN_6815 = {{24'd0}, _T_25744};
  assign _T_65799 = _GEN_6815 << 24;
  assign _GEN_6816 = {{8'd0}, _T_65763};
  assign _T_65803 = _GEN_6816 | _T_65799;
  assign _GEN_6817 = {{8'd0}, _T_25204};
  assign _T_65879 = _GEN_6817 << 8;
  assign _GEN_6818 = {{8'd0}, _T_25202};
  assign _T_65883 = _GEN_6818 | _T_65879;
  assign _GEN_6819 = {{16'd0}, _T_25206};
  assign _T_65919 = _GEN_6819 << 16;
  assign _GEN_6820 = {{8'd0}, _T_65883};
  assign _T_65923 = _GEN_6820 | _T_65919;
  assign _GEN_6821 = {{24'd0}, _T_25208};
  assign _T_65959 = _GEN_6821 << 24;
  assign _GEN_6822 = {{8'd0}, _T_65923};
  assign _T_65963 = _GEN_6822 | _T_65959;
  assign _GEN_6823 = {{8'd0}, _T_25148};
  assign _T_66039 = _GEN_6823 << 8;
  assign _GEN_6824 = {{8'd0}, _T_25146};
  assign _T_66043 = _GEN_6824 | _T_66039;
  assign _GEN_6825 = {{16'd0}, _T_25150};
  assign _T_66079 = _GEN_6825 << 16;
  assign _GEN_6826 = {{8'd0}, _T_66043};
  assign _T_66083 = _GEN_6826 | _T_66079;
  assign _GEN_6827 = {{24'd0}, _T_25152};
  assign _T_66119 = _GEN_6827 << 24;
  assign _GEN_6828 = {{8'd0}, _T_66083};
  assign _T_66123 = _GEN_6828 | _T_66119;
  assign _GEN_6829 = {{8'd0}, _T_25484};
  assign _T_66199 = _GEN_6829 << 8;
  assign _GEN_6830 = {{8'd0}, _T_25482};
  assign _T_66203 = _GEN_6830 | _T_66199;
  assign _GEN_6831 = {{16'd0}, _T_25486};
  assign _T_66239 = _GEN_6831 << 16;
  assign _GEN_6832 = {{8'd0}, _T_66203};
  assign _T_66243 = _GEN_6832 | _T_66239;
  assign _GEN_6833 = {{24'd0}, _T_25488};
  assign _T_66279 = _GEN_6833 << 24;
  assign _GEN_6834 = {{8'd0}, _T_66243};
  assign _T_66283 = _GEN_6834 | _T_66279;
  assign _GEN_6835 = {{8'd0}, _T_25620};
  assign _T_66359 = _GEN_6835 << 8;
  assign _GEN_6836 = {{8'd0}, _T_25618};
  assign _T_66363 = _GEN_6836 | _T_66359;
  assign _GEN_6837 = {{16'd0}, _T_25622};
  assign _T_66399 = _GEN_6837 << 16;
  assign _GEN_6838 = {{8'd0}, _T_66363};
  assign _T_66403 = _GEN_6838 | _T_66399;
  assign _GEN_6839 = {{24'd0}, _T_25624};
  assign _T_66439 = _GEN_6839 << 24;
  assign _GEN_6840 = {{8'd0}, _T_66403};
  assign _T_66443 = _GEN_6840 | _T_66439;
  assign _GEN_6841 = {{8'd0}, _T_25108};
  assign _T_66519 = _GEN_6841 << 8;
  assign _GEN_6842 = {{8'd0}, _T_25106};
  assign _T_66523 = _GEN_6842 | _T_66519;
  assign _GEN_6843 = {{16'd0}, _T_25110};
  assign _T_66559 = _GEN_6843 << 16;
  assign _GEN_6844 = {{8'd0}, _T_66523};
  assign _T_66563 = _GEN_6844 | _T_66559;
  assign _GEN_6845 = {{24'd0}, _T_25112};
  assign _T_66599 = _GEN_6845 << 24;
  assign _GEN_6846 = {{8'd0}, _T_66563};
  assign _T_66603 = _GEN_6846 | _T_66599;
  assign _GEN_6847 = {{8'd0}, _T_24692};
  assign _T_66839 = _GEN_6847 << 8;
  assign _GEN_6848 = {{8'd0}, _T_24690};
  assign _T_66843 = _GEN_6848 | _T_66839;
  assign _GEN_6849 = {{16'd0}, _T_24694};
  assign _T_66879 = _GEN_6849 << 16;
  assign _GEN_6850 = {{8'd0}, _T_66843};
  assign _T_66883 = _GEN_6850 | _T_66879;
  assign _GEN_6851 = {{24'd0}, _T_24696};
  assign _T_66919 = _GEN_6851 << 24;
  assign _GEN_6852 = {{8'd0}, _T_66883};
  assign _T_66923 = _GEN_6852 | _T_66919;
  assign _T_66943 = _T_99434 & _T_35050;
  assign _GEN_2486 = _T_66943 ? _T_35064 : _GEN_325;
  assign _T_66983 = _T_99434 & _T_35090;
  assign _GEN_2487 = _T_66983 ? _T_35104 : _GEN_326;
  assign _T_67023 = _T_99434 & _T_35130;
  assign _GEN_2488 = _T_67023 ? _T_35144 : _GEN_327;
  assign _T_67063 = _T_99434 & _T_35170;
  assign _GEN_2489 = _T_67063 ? _T_35184 : _GEN_328;
  assign _GEN_6859 = {{8'd0}, _T_25596};
  assign _T_67159 = _GEN_6859 << 8;
  assign _GEN_6860 = {{8'd0}, _T_25594};
  assign _T_67163 = _GEN_6860 | _T_67159;
  assign _GEN_6861 = {{16'd0}, _T_25598};
  assign _T_67199 = _GEN_6861 << 16;
  assign _GEN_6862 = {{8'd0}, _T_67163};
  assign _T_67203 = _GEN_6862 | _T_67199;
  assign _GEN_6863 = {{24'd0}, _T_25600};
  assign _T_67239 = _GEN_6863 << 24;
  assign _GEN_6864 = {{8'd0}, _T_67203};
  assign _T_67243 = _GEN_6864 | _T_67239;
  assign _GEN_6865 = {{8'd0}, _T_24436};
  assign _T_67479 = _GEN_6865 << 8;
  assign _GEN_6866 = {{8'd0}, _T_24434};
  assign _T_67483 = _GEN_6866 | _T_67479;
  assign _GEN_6867 = {{16'd0}, _T_24438};
  assign _T_67519 = _GEN_6867 << 16;
  assign _GEN_6868 = {{8'd0}, _T_67483};
  assign _T_67523 = _GEN_6868 | _T_67519;
  assign _GEN_6869 = {{24'd0}, _T_24440};
  assign _T_67559 = _GEN_6869 << 24;
  assign _GEN_6870 = {{8'd0}, _T_67523};
  assign _T_67563 = _GEN_6870 | _T_67559;
  assign _GEN_6871 = {{8'd0}, _T_24540};
  assign _T_67639 = _GEN_6871 << 8;
  assign _GEN_6872 = {{8'd0}, _T_24538};
  assign _T_67643 = _GEN_6872 | _T_67639;
  assign _GEN_6873 = {{16'd0}, _T_24542};
  assign _T_67679 = _GEN_6873 << 16;
  assign _GEN_6874 = {{8'd0}, _T_67643};
  assign _T_67683 = _GEN_6874 | _T_67679;
  assign _GEN_6875 = {{24'd0}, _T_24544};
  assign _T_67719 = _GEN_6875 << 24;
  assign _GEN_6876 = {{8'd0}, _T_67683};
  assign _T_67723 = _GEN_6876 | _T_67719;
  assign _GEN_6877 = {{8'd0}, _T_25364};
  assign _T_67799 = _GEN_6877 << 8;
  assign _GEN_6878 = {{8'd0}, _T_25362};
  assign _T_67803 = _GEN_6878 | _T_67799;
  assign _GEN_6879 = {{16'd0}, _T_25366};
  assign _T_67839 = _GEN_6879 << 16;
  assign _GEN_6880 = {{8'd0}, _T_67803};
  assign _T_67843 = _GEN_6880 | _T_67839;
  assign _GEN_6881 = {{24'd0}, _T_25368};
  assign _T_67879 = _GEN_6881 << 24;
  assign _GEN_6882 = {{8'd0}, _T_67843};
  assign _T_67883 = _GEN_6882 | _T_67879;
  assign _GEN_6883 = {{8'd0}, _T_24060};
  assign _T_68119 = _GEN_6883 << 8;
  assign _GEN_6884 = {{8'd0}, _T_24058};
  assign _T_68123 = _GEN_6884 | _T_68119;
  assign _GEN_6885 = {{16'd0}, _T_24062};
  assign _T_68159 = _GEN_6885 << 16;
  assign _GEN_6886 = {{8'd0}, _T_68123};
  assign _T_68163 = _GEN_6886 | _T_68159;
  assign _GEN_6887 = {{24'd0}, _T_24064};
  assign _T_68199 = _GEN_6887 << 24;
  assign _GEN_6888 = {{8'd0}, _T_68163};
  assign _T_68203 = _GEN_6888 | _T_68199;
  assign _GEN_6889 = {{8'd0}, _T_23956};
  assign _T_68279 = _GEN_6889 << 8;
  assign _GEN_6890 = {{8'd0}, _T_23954};
  assign _T_68283 = _GEN_6890 | _T_68279;
  assign _GEN_6891 = {{16'd0}, _T_23958};
  assign _T_68319 = _GEN_6891 << 16;
  assign _GEN_6892 = {{8'd0}, _T_68283};
  assign _T_68323 = _GEN_6892 | _T_68319;
  assign _GEN_6893 = {{24'd0}, _T_23960};
  assign _T_68359 = _GEN_6893 << 24;
  assign _GEN_6894 = {{8'd0}, _T_68323};
  assign _T_68363 = _GEN_6894 | _T_68359;
  assign _GEN_6895 = {{8'd0}, _T_25012};
  assign _T_68439 = _GEN_6895 << 8;
  assign _GEN_6896 = {{8'd0}, _T_25010};
  assign _T_68443 = _GEN_6896 | _T_68439;
  assign _GEN_6897 = {{16'd0}, _T_25014};
  assign _T_68479 = _GEN_6897 << 16;
  assign _GEN_6898 = {{8'd0}, _T_68443};
  assign _T_68483 = _GEN_6898 | _T_68479;
  assign _GEN_6899 = {{24'd0}, _T_25016};
  assign _T_68519 = _GEN_6899 << 24;
  assign _GEN_6900 = {{8'd0}, _T_68483};
  assign _T_68523 = _GEN_6900 | _T_68519;
  assign _GEN_6901 = {{8'd0}, _T_24316};
  assign _T_68599 = _GEN_6901 << 8;
  assign _GEN_6902 = {{8'd0}, _T_24314};
  assign _T_68603 = _GEN_6902 | _T_68599;
  assign _GEN_6903 = {{16'd0}, _T_24318};
  assign _T_68639 = _GEN_6903 << 16;
  assign _GEN_6904 = {{8'd0}, _T_68603};
  assign _T_68643 = _GEN_6904 | _T_68639;
  assign _GEN_6905 = {{24'd0}, _T_24320};
  assign _T_68679 = _GEN_6905 << 24;
  assign _GEN_6906 = {{8'd0}, _T_68643};
  assign _T_68683 = _GEN_6906 | _T_68679;
  assign _GEN_6907 = {{8'd0}, _T_24972};
  assign _T_68759 = _GEN_6907 << 8;
  assign _GEN_6908 = {{8'd0}, _T_24970};
  assign _T_68763 = _GEN_6908 | _T_68759;
  assign _GEN_6909 = {{16'd0}, _T_24974};
  assign _T_68799 = _GEN_6909 << 16;
  assign _GEN_6910 = {{8'd0}, _T_68763};
  assign _T_68803 = _GEN_6910 | _T_68799;
  assign _GEN_6911 = {{24'd0}, _T_24976};
  assign _T_68839 = _GEN_6911 << 24;
  assign _GEN_6912 = {{8'd0}, _T_68803};
  assign _T_68843 = _GEN_6912 | _T_68839;
  assign _GEN_6913 = {{8'd0}, _T_23804};
  assign _T_68919 = _GEN_6913 << 8;
  assign _GEN_6914 = {{8'd0}, _T_23802};
  assign _T_68923 = _GEN_6914 | _T_68919;
  assign _GEN_6915 = {{16'd0}, _T_23806};
  assign _T_68959 = _GEN_6915 << 16;
  assign _GEN_6916 = {{8'd0}, _T_68923};
  assign _T_68963 = _GEN_6916 | _T_68959;
  assign _GEN_6917 = {{24'd0}, _T_23808};
  assign _T_68999 = _GEN_6917 << 24;
  assign _GEN_6918 = {{8'd0}, _T_68963};
  assign _T_69003 = _GEN_6918 | _T_68999;
  assign _GEN_6919 = {{8'd0}, _T_24180};
  assign _T_69079 = _GEN_6919 << 8;
  assign _GEN_6920 = {{8'd0}, _T_24178};
  assign _T_69083 = _GEN_6920 | _T_69079;
  assign _GEN_6921 = {{16'd0}, _T_24182};
  assign _T_69119 = _GEN_6921 << 16;
  assign _GEN_6922 = {{8'd0}, _T_69083};
  assign _T_69123 = _GEN_6922 | _T_69119;
  assign _GEN_6923 = {{24'd0}, _T_24184};
  assign _T_69159 = _GEN_6923 << 24;
  assign _GEN_6924 = {{8'd0}, _T_69123};
  assign _T_69163 = _GEN_6924 | _T_69159;
  assign _T_69183 = _T_98298 & _T_50170;
  assign _GEN_6925 = {{8'd0}, _T_24348};
  assign _T_69279 = _GEN_6925 << 8;
  assign _GEN_6926 = {{8'd0}, _T_24346};
  assign _T_69283 = _GEN_6926 | _T_69279;
  assign _GEN_6927 = {{16'd0}, _T_24350};
  assign _T_69319 = _GEN_6927 << 16;
  assign _GEN_6928 = {{8'd0}, _T_69283};
  assign _T_69323 = _GEN_6928 | _T_69319;
  assign _GEN_6929 = {{24'd0}, _T_24352};
  assign _T_69359 = _GEN_6929 << 24;
  assign _GEN_6930 = {{8'd0}, _T_69323};
  assign _T_69363 = _GEN_6930 | _T_69359;
  assign _GEN_6931 = {{8'd0}, _T_25228};
  assign _T_69439 = _GEN_6931 << 8;
  assign _GEN_6932 = {{8'd0}, _T_25226};
  assign _T_69443 = _GEN_6932 | _T_69439;
  assign _GEN_6933 = {{16'd0}, _T_25230};
  assign _T_69479 = _GEN_6933 << 16;
  assign _GEN_6934 = {{8'd0}, _T_69443};
  assign _T_69483 = _GEN_6934 | _T_69479;
  assign _GEN_6935 = {{24'd0}, _T_25232};
  assign _T_69519 = _GEN_6935 << 24;
  assign _GEN_6936 = {{8'd0}, _T_69483};
  assign _T_69523 = _GEN_6936 | _T_69519;
  assign _GEN_6937 = {{8'd0}, _T_24660};
  assign _T_69599 = _GEN_6937 << 8;
  assign _GEN_6938 = {{8'd0}, _T_24658};
  assign _T_69603 = _GEN_6938 | _T_69599;
  assign _GEN_6939 = {{16'd0}, _T_24662};
  assign _T_69639 = _GEN_6939 << 16;
  assign _GEN_6940 = {{8'd0}, _T_69603};
  assign _T_69643 = _GEN_6940 | _T_69639;
  assign _GEN_6941 = {{24'd0}, _T_24664};
  assign _T_69679 = _GEN_6941 << 24;
  assign _GEN_6942 = {{8'd0}, _T_69643};
  assign _T_69683 = _GEN_6942 | _T_69679;
  assign _GEN_6943 = {{8'd0}, _T_25716};
  assign _T_69759 = _GEN_6943 << 8;
  assign _GEN_6944 = {{8'd0}, _T_25714};
  assign _T_69763 = _GEN_6944 | _T_69759;
  assign _GEN_6945 = {{16'd0}, _T_25718};
  assign _T_69799 = _GEN_6945 << 16;
  assign _GEN_6946 = {{8'd0}, _T_69763};
  assign _T_69803 = _GEN_6946 | _T_69799;
  assign _GEN_6947 = {{24'd0}, _T_25720};
  assign _T_69839 = _GEN_6947 << 24;
  assign _GEN_6948 = {{8'd0}, _T_69803};
  assign _T_69843 = _GEN_6948 | _T_69839;
  assign _GEN_6949 = {{8'd0}, _T_25404};
  assign _T_69919 = _GEN_6949 << 8;
  assign _GEN_6950 = {{8'd0}, _T_25402};
  assign _T_69923 = _GEN_6950 | _T_69919;
  assign _GEN_6951 = {{16'd0}, _T_25406};
  assign _T_69959 = _GEN_6951 << 16;
  assign _GEN_6952 = {{8'd0}, _T_69923};
  assign _T_69963 = _GEN_6952 | _T_69959;
  assign _GEN_6953 = {{24'd0}, _T_25408};
  assign _T_69999 = _GEN_6953 << 24;
  assign _GEN_6954 = {{8'd0}, _T_69963};
  assign _T_70003 = _GEN_6954 | _T_69999;
  assign _GEN_6955 = {{8'd0}, _T_24404};
  assign _T_70079 = _GEN_6955 << 8;
  assign _GEN_6956 = {{8'd0}, _T_24402};
  assign _T_70083 = _GEN_6956 | _T_70079;
  assign _GEN_6957 = {{16'd0}, _T_24406};
  assign _T_70119 = _GEN_6957 << 16;
  assign _GEN_6958 = {{8'd0}, _T_70083};
  assign _T_70123 = _GEN_6958 | _T_70119;
  assign _GEN_6959 = {{24'd0}, _T_24408};
  assign _T_70159 = _GEN_6959 << 24;
  assign _GEN_6960 = {{8'd0}, _T_70123};
  assign _T_70163 = _GEN_6960 | _T_70159;
  assign _GEN_6961 = {{8'd0}, _T_25460};
  assign _T_70239 = _GEN_6961 << 8;
  assign _GEN_6962 = {{8'd0}, _T_25458};
  assign _T_70243 = _GEN_6962 | _T_70239;
  assign _GEN_6963 = {{16'd0}, _T_25462};
  assign _T_70279 = _GEN_6963 << 16;
  assign _GEN_6964 = {{8'd0}, _T_70243};
  assign _T_70283 = _GEN_6964 | _T_70279;
  assign _GEN_6965 = {{24'd0}, _T_25464};
  assign _T_70319 = _GEN_6965 << 24;
  assign _GEN_6966 = {{8'd0}, _T_70283};
  assign _T_70323 = _GEN_6966 | _T_70319;
  assign _GEN_6967 = {{8'd0}, _T_24572};
  assign _T_70399 = _GEN_6967 << 8;
  assign _GEN_6968 = {{8'd0}, _T_24570};
  assign _T_70403 = _GEN_6968 | _T_70399;
  assign _GEN_6969 = {{16'd0}, _T_24574};
  assign _T_70439 = _GEN_6969 << 16;
  assign _GEN_6970 = {{8'd0}, _T_70403};
  assign _T_70443 = _GEN_6970 | _T_70439;
  assign _GEN_6971 = {{24'd0}, _T_24576};
  assign _T_70479 = _GEN_6971 << 24;
  assign _GEN_6972 = {{8'd0}, _T_70443};
  assign _T_70483 = _GEN_6972 | _T_70479;
  assign _GEN_6973 = {{8'd0}, _T_24388};
  assign _T_70559 = _GEN_6973 << 8;
  assign _GEN_6974 = {{8'd0}, _T_24386};
  assign _T_70563 = _GEN_6974 | _T_70559;
  assign _GEN_6975 = {{16'd0}, _T_24390};
  assign _T_70599 = _GEN_6975 << 16;
  assign _GEN_6976 = {{8'd0}, _T_70563};
  assign _T_70603 = _GEN_6976 | _T_70599;
  assign _GEN_6977 = {{24'd0}, _T_24392};
  assign _T_70639 = _GEN_6977 << 24;
  assign _GEN_6978 = {{8'd0}, _T_70603};
  assign _T_70643 = _GEN_6978 | _T_70639;
  assign _GEN_6979 = {{8'd0}, _T_24788};
  assign _T_70719 = _GEN_6979 << 8;
  assign _GEN_6980 = {{8'd0}, _T_24786};
  assign _T_70723 = _GEN_6980 | _T_70719;
  assign _GEN_6981 = {{16'd0}, _T_24790};
  assign _T_70759 = _GEN_6981 << 16;
  assign _GEN_6982 = {{8'd0}, _T_70723};
  assign _T_70763 = _GEN_6982 | _T_70759;
  assign _GEN_6983 = {{24'd0}, _T_24792};
  assign _T_70799 = _GEN_6983 << 24;
  assign _GEN_6984 = {{8'd0}, _T_70763};
  assign _T_70803 = _GEN_6984 | _T_70799;
  assign _GEN_6985 = {{8'd0}, _T_24212};
  assign _T_70879 = _GEN_6985 << 8;
  assign _GEN_6986 = {{8'd0}, _T_24210};
  assign _T_70883 = _GEN_6986 | _T_70879;
  assign _GEN_6987 = {{16'd0}, _T_24214};
  assign _T_70919 = _GEN_6987 << 16;
  assign _GEN_6988 = {{8'd0}, _T_70883};
  assign _T_70923 = _GEN_6988 | _T_70919;
  assign _GEN_6989 = {{24'd0}, _T_24216};
  assign _T_70959 = _GEN_6989 << 24;
  assign _GEN_6990 = {{8'd0}, _T_70923};
  assign _T_70963 = _GEN_6990 | _T_70959;
  assign _GEN_6991 = {{8'd0}, _T_25268};
  assign _T_71039 = _GEN_6991 << 8;
  assign _GEN_6992 = {{8'd0}, _T_25266};
  assign _T_71043 = _GEN_6992 | _T_71039;
  assign _GEN_6993 = {{16'd0}, _T_25270};
  assign _T_71079 = _GEN_6993 << 16;
  assign _GEN_6994 = {{8'd0}, _T_71043};
  assign _T_71083 = _GEN_6994 | _T_71079;
  assign _GEN_6995 = {{24'd0}, _T_25272};
  assign _T_71119 = _GEN_6995 << 24;
  assign _GEN_6996 = {{8'd0}, _T_71083};
  assign _T_71123 = _GEN_6996 | _T_71119;
  assign _GEN_6997 = {{8'd0}, _T_25676};
  assign _T_71199 = _GEN_6997 << 8;
  assign _GEN_6998 = {{8'd0}, _T_25674};
  assign _T_71203 = _GEN_6998 | _T_71199;
  assign _GEN_6999 = {{16'd0}, _T_25678};
  assign _T_71239 = _GEN_6999 << 16;
  assign _GEN_7000 = {{8'd0}, _T_71203};
  assign _T_71243 = _GEN_7000 | _T_71239;
  assign _GEN_7001 = {{24'd0}, _T_25680};
  assign _T_71279 = _GEN_7001 << 24;
  assign _GEN_7002 = {{8'd0}, _T_71243};
  assign _T_71283 = _GEN_7002 | _T_71279;
  assign _GEN_7003 = {{8'd0}, _T_25420};
  assign _T_71359 = _GEN_7003 << 8;
  assign _GEN_7004 = {{8'd0}, _T_25418};
  assign _T_71363 = _GEN_7004 | _T_71359;
  assign _GEN_7005 = {{16'd0}, _T_25422};
  assign _T_71399 = _GEN_7005 << 16;
  assign _GEN_7006 = {{8'd0}, _T_71363};
  assign _T_71403 = _GEN_7006 | _T_71399;
  assign _GEN_7007 = {{24'd0}, _T_25424};
  assign _T_71439 = _GEN_7007 << 24;
  assign _GEN_7008 = {{8'd0}, _T_71403};
  assign _T_71443 = _GEN_7008 | _T_71439;
  assign _GEN_7009 = {{8'd0}, _T_25300};
  assign _T_71519 = _GEN_7009 << 8;
  assign _GEN_7010 = {{8'd0}, _T_25298};
  assign _T_71523 = _GEN_7010 | _T_71519;
  assign _GEN_7011 = {{16'd0}, _T_25302};
  assign _T_71559 = _GEN_7011 << 16;
  assign _GEN_7012 = {{8'd0}, _T_71523};
  assign _T_71563 = _GEN_7012 | _T_71559;
  assign _GEN_7013 = {{24'd0}, _T_25304};
  assign _T_71599 = _GEN_7013 << 24;
  assign _GEN_7014 = {{8'd0}, _T_71563};
  assign _T_71603 = _GEN_7014 | _T_71599;
  assign _GEN_7015 = {{8'd0}, _T_24604};
  assign _T_71679 = _GEN_7015 << 8;
  assign _GEN_7016 = {{8'd0}, _T_24602};
  assign _T_71683 = _GEN_7016 | _T_71679;
  assign _GEN_7017 = {{16'd0}, _T_24606};
  assign _T_71719 = _GEN_7017 << 16;
  assign _GEN_7018 = {{8'd0}, _T_71683};
  assign _T_71723 = _GEN_7018 | _T_71719;
  assign _GEN_7019 = {{24'd0}, _T_24608};
  assign _T_71759 = _GEN_7019 << 24;
  assign _GEN_7020 = {{8'd0}, _T_71723};
  assign _T_71763 = _GEN_7020 | _T_71759;
  assign _GEN_7021 = {{8'd0}, _T_25556};
  assign _T_71839 = _GEN_7021 << 8;
  assign _GEN_7022 = {{8'd0}, _T_25554};
  assign _T_71843 = _GEN_7022 | _T_71839;
  assign _GEN_7023 = {{16'd0}, _T_25558};
  assign _T_71879 = _GEN_7023 << 16;
  assign _GEN_7024 = {{8'd0}, _T_71843};
  assign _T_71883 = _GEN_7024 | _T_71879;
  assign _GEN_7025 = {{24'd0}, _T_25560};
  assign _T_71919 = _GEN_7025 << 24;
  assign _GEN_7026 = {{8'd0}, _T_71883};
  assign _T_71923 = _GEN_7026 | _T_71919;
  assign _GEN_7027 = {{8'd0}, _T_25660};
  assign _T_72159 = _GEN_7027 << 8;
  assign _GEN_7028 = {{8'd0}, _T_25658};
  assign _T_72163 = _GEN_7028 | _T_72159;
  assign _GEN_7029 = {{16'd0}, _T_25662};
  assign _T_72199 = _GEN_7029 << 16;
  assign _GEN_7030 = {{8'd0}, _T_72163};
  assign _T_72203 = _GEN_7030 | _T_72199;
  assign _GEN_7031 = {{24'd0}, _T_25664};
  assign _T_72239 = _GEN_7031 << 24;
  assign _GEN_7032 = {{8'd0}, _T_72203};
  assign _T_72243 = _GEN_7032 | _T_72239;
  assign _T_72263 = _T_99506 & _T_35050;
  assign _GEN_2491 = _T_72263 ? _T_35064 : _GEN_361;
  assign _T_72303 = _T_99506 & _T_35090;
  assign _GEN_2492 = _T_72303 ? _T_35104 : _GEN_362;
  assign _T_72343 = _T_99506 & _T_35130;
  assign _GEN_2493 = _T_72343 ? _T_35144 : _GEN_363;
  assign _T_72383 = _T_99506 & _T_35170;
  assign _GEN_2494 = _T_72383 ? _T_35184 : _GEN_364;
  assign _GEN_7039 = {{8'd0}, _T_24644};
  assign _T_72479 = _GEN_7039 << 8;
  assign _GEN_7040 = {{8'd0}, _T_24642};
  assign _T_72483 = _GEN_7040 | _T_72479;
  assign _GEN_7041 = {{16'd0}, _T_24646};
  assign _T_72519 = _GEN_7041 << 16;
  assign _GEN_7042 = {{8'd0}, _T_72483};
  assign _T_72523 = _GEN_7042 | _T_72519;
  assign _GEN_7043 = {{24'd0}, _T_24648};
  assign _T_72559 = _GEN_7043 << 24;
  assign _GEN_7044 = {{8'd0}, _T_72523};
  assign _T_72563 = _GEN_7044 | _T_72559;
  assign _GEN_7045 = {{8'd0}, _T_24252};
  assign _T_72799 = _GEN_7045 << 8;
  assign _GEN_7046 = {{8'd0}, _T_24250};
  assign _T_72803 = _GEN_7046 | _T_72799;
  assign _GEN_7047 = {{16'd0}, _T_24254};
  assign _T_72839 = _GEN_7047 << 16;
  assign _GEN_7048 = {{8'd0}, _T_72803};
  assign _T_72843 = _GEN_7048 | _T_72839;
  assign _GEN_7049 = {{24'd0}, _T_24256};
  assign _T_72879 = _GEN_7049 << 24;
  assign _GEN_7050 = {{8'd0}, _T_72843};
  assign _T_72883 = _GEN_7050 | _T_72879;
  assign _GEN_7051 = {{8'd0}, _T_24132};
  assign _T_72959 = _GEN_7051 << 8;
  assign _GEN_7052 = {{8'd0}, _T_24130};
  assign _T_72963 = _GEN_7052 | _T_72959;
  assign _GEN_7053 = {{16'd0}, _T_24134};
  assign _T_72999 = _GEN_7053 << 16;
  assign _GEN_7054 = {{8'd0}, _T_72963};
  assign _T_73003 = _GEN_7054 | _T_72999;
  assign _GEN_7055 = {{24'd0}, _T_24136};
  assign _T_73039 = _GEN_7055 << 24;
  assign _GEN_7056 = {{8'd0}, _T_73003};
  assign _T_73043 = _GEN_7056 | _T_73039;
  assign _GEN_7057 = {{8'd0}, _T_23764};
  assign _T_73119 = _GEN_7057 << 8;
  assign _GEN_7058 = {{8'd0}, _T_23762};
  assign _T_73123 = _GEN_7058 | _T_73119;
  assign _GEN_7059 = {{16'd0}, _T_23766};
  assign _T_73159 = _GEN_7059 << 16;
  assign _GEN_7060 = {{8'd0}, _T_73123};
  assign _T_73163 = _GEN_7060 | _T_73159;
  assign _GEN_7061 = {{24'd0}, _T_23768};
  assign _T_73199 = _GEN_7061 << 24;
  assign _GEN_7062 = {{8'd0}, _T_73163};
  assign _T_73203 = _GEN_7062 | _T_73199;
  assign _GEN_7063 = {{8'd0}, _T_24508};
  assign _T_73279 = _GEN_7063 << 8;
  assign _GEN_7064 = {{8'd0}, _T_24506};
  assign _T_73283 = _GEN_7064 | _T_73279;
  assign _GEN_7065 = {{16'd0}, _T_24510};
  assign _T_73319 = _GEN_7065 << 16;
  assign _GEN_7066 = {{8'd0}, _T_73283};
  assign _T_73323 = _GEN_7066 | _T_73319;
  assign _GEN_7067 = {{24'd0}, _T_24512};
  assign _T_73359 = _GEN_7067 << 24;
  assign _GEN_7068 = {{8'd0}, _T_73323};
  assign _T_73363 = _GEN_7068 | _T_73359;
  assign _GEN_7069 = {{8'd0}, _T_24820};
  assign _T_73439 = _GEN_7069 << 8;
  assign _GEN_7070 = {{8'd0}, _T_24818};
  assign _T_73443 = _GEN_7070 | _T_73439;
  assign _GEN_7071 = {{16'd0}, _T_24822};
  assign _T_73479 = _GEN_7071 << 16;
  assign _GEN_7072 = {{8'd0}, _T_73443};
  assign _T_73483 = _GEN_7072 | _T_73479;
  assign _GEN_7073 = {{24'd0}, _T_24824};
  assign _T_73519 = _GEN_7073 << 24;
  assign _GEN_7074 = {{8'd0}, _T_73483};
  assign _T_73523 = _GEN_7074 | _T_73519;
  assign _GEN_7075 = {{8'd0}, _T_24908};
  assign _T_73599 = _GEN_7075 << 8;
  assign _GEN_7076 = {{8'd0}, _T_24906};
  assign _T_73603 = _GEN_7076 | _T_73599;
  assign _GEN_7077 = {{16'd0}, _T_24910};
  assign _T_73639 = _GEN_7077 << 16;
  assign _GEN_7078 = {{8'd0}, _T_73603};
  assign _T_73643 = _GEN_7078 | _T_73639;
  assign _GEN_7079 = {{24'd0}, _T_24912};
  assign _T_73679 = _GEN_7079 << 24;
  assign _GEN_7080 = {{8'd0}, _T_73643};
  assign _T_73683 = _GEN_7080 | _T_73679;
  assign _GEN_7081 = {{8'd0}, _T_25044};
  assign _T_73759 = _GEN_7081 << 8;
  assign _GEN_7082 = {{8'd0}, _T_25042};
  assign _T_73763 = _GEN_7082 | _T_73759;
  assign _GEN_7083 = {{16'd0}, _T_25046};
  assign _T_73799 = _GEN_7083 << 16;
  assign _GEN_7084 = {{8'd0}, _T_73763};
  assign _T_73803 = _GEN_7084 | _T_73799;
  assign _GEN_7085 = {{24'd0}, _T_25048};
  assign _T_73839 = _GEN_7085 << 24;
  assign _GEN_7086 = {{8'd0}, _T_73803};
  assign _T_73843 = _GEN_7086 | _T_73839;
  assign _GEN_7087 = {{8'd0}, _T_24020};
  assign _T_73919 = _GEN_7087 << 8;
  assign _GEN_7088 = {{8'd0}, _T_24018};
  assign _T_73923 = _GEN_7088 | _T_73919;
  assign _GEN_7089 = {{16'd0}, _T_24022};
  assign _T_73959 = _GEN_7089 << 16;
  assign _GEN_7090 = {{8'd0}, _T_73923};
  assign _T_73963 = _GEN_7090 | _T_73959;
  assign _GEN_7091 = {{24'd0}, _T_24024};
  assign _T_73999 = _GEN_7091 << 24;
  assign _GEN_7092 = {{8'd0}, _T_73963};
  assign _T_74003 = _GEN_7092 | _T_73999;
  assign _GEN_7093 = {{8'd0}, _T_24724};
  assign _T_74079 = _GEN_7093 << 8;
  assign _GEN_7094 = {{8'd0}, _T_24722};
  assign _T_74083 = _GEN_7094 | _T_74079;
  assign _GEN_7095 = {{16'd0}, _T_24726};
  assign _T_74119 = _GEN_7095 << 16;
  assign _GEN_7096 = {{8'd0}, _T_74083};
  assign _T_74123 = _GEN_7096 | _T_74119;
  assign _GEN_7097 = {{24'd0}, _T_24728};
  assign _T_74159 = _GEN_7097 << 24;
  assign _GEN_7098 = {{8'd0}, _T_74123};
  assign _T_74163 = _GEN_7098 | _T_74159;
  assign _GEN_7099 = {{8'd0}, _T_25164};
  assign _T_74239 = _GEN_7099 << 8;
  assign _GEN_7100 = {{8'd0}, _T_25162};
  assign _T_74243 = _GEN_7100 | _T_74239;
  assign _GEN_7101 = {{16'd0}, _T_25166};
  assign _T_74279 = _GEN_7101 << 16;
  assign _GEN_7102 = {{8'd0}, _T_74243};
  assign _T_74283 = _GEN_7102 | _T_74279;
  assign _GEN_7103 = {{24'd0}, _T_25168};
  assign _T_74319 = _GEN_7103 << 24;
  assign _GEN_7104 = {{8'd0}, _T_74283};
  assign _T_74323 = _GEN_7104 | _T_74319;
  assign _GEN_7105 = {{8'd0}, _T_25780};
  assign _T_74399 = _GEN_7105 << 8;
  assign _GEN_7106 = {{8'd0}, _T_25778};
  assign _T_74403 = _GEN_7106 | _T_74399;
  assign _GEN_7107 = {{16'd0}, _T_25782};
  assign _T_74439 = _GEN_7107 << 16;
  assign _GEN_7108 = {{8'd0}, _T_74403};
  assign _T_74443 = _GEN_7108 | _T_74439;
  assign _GEN_7109 = {{24'd0}, _T_25784};
  assign _T_74479 = _GEN_7109 << 24;
  assign _GEN_7110 = {{8'd0}, _T_74443};
  assign _T_74483 = _GEN_7110 | _T_74479;
  assign _GEN_7111 = {{8'd0}, _T_25524};
  assign _T_74599 = _GEN_7111 << 8;
  assign _GEN_7112 = {{8'd0}, _T_25522};
  assign _T_74603 = _GEN_7112 | _T_74599;
  assign _GEN_7113 = {{16'd0}, _T_25526};
  assign _T_74639 = _GEN_7113 << 16;
  assign _GEN_7114 = {{8'd0}, _T_74603};
  assign _T_74643 = _GEN_7114 | _T_74639;
  assign _GEN_7115 = {{24'd0}, _T_25528};
  assign _T_74679 = _GEN_7115 << 24;
  assign _GEN_7116 = {{8'd0}, _T_74643};
  assign _T_74683 = _GEN_7116 | _T_74679;
  assign _GEN_7117 = {{8'd0}, _T_23876};
  assign _T_74759 = _GEN_7117 << 8;
  assign _GEN_7118 = {{8'd0}, _T_23874};
  assign _T_74763 = _GEN_7118 | _T_74759;
  assign _GEN_7119 = {{16'd0}, _T_23878};
  assign _T_74799 = _GEN_7119 << 16;
  assign _GEN_7120 = {{8'd0}, _T_74763};
  assign _T_74803 = _GEN_7120 | _T_74799;
  assign _GEN_7121 = {{24'd0}, _T_23880};
  assign _T_74839 = _GEN_7121 << 24;
  assign _GEN_7122 = {{8'd0}, _T_74803};
  assign _T_74843 = _GEN_7122 | _T_74839;
  assign _GEN_7123 = {{8'd0}, _T_24764};
  assign _T_74919 = _GEN_7123 << 8;
  assign _GEN_7124 = {{8'd0}, _T_24762};
  assign _T_74923 = _GEN_7124 | _T_74919;
  assign _GEN_7125 = {{16'd0}, _T_24766};
  assign _T_74959 = _GEN_7125 << 16;
  assign _GEN_7126 = {{8'd0}, _T_74923};
  assign _T_74963 = _GEN_7126 | _T_74959;
  assign _GEN_7127 = {{24'd0}, _T_24768};
  assign _T_74999 = _GEN_7127 << 24;
  assign _GEN_7128 = {{8'd0}, _T_74963};
  assign _T_75003 = _GEN_7128 | _T_74999;
  assign _GEN_7129 = {{8'd0}, _T_24468};
  assign _T_75079 = _GEN_7129 << 8;
  assign _GEN_7130 = {{8'd0}, _T_24466};
  assign _T_75083 = _GEN_7130 | _T_75079;
  assign _GEN_7131 = {{16'd0}, _T_24470};
  assign _T_75119 = _GEN_7131 << 16;
  assign _GEN_7132 = {{8'd0}, _T_75083};
  assign _T_75123 = _GEN_7132 | _T_75119;
  assign _GEN_7133 = {{24'd0}, _T_24472};
  assign _T_75159 = _GEN_7133 << 24;
  assign _GEN_7134 = {{8'd0}, _T_75123};
  assign _T_75163 = _GEN_7134 | _T_75159;
  assign _T_75183 = _T_99474 & _T_35050;
  assign _GEN_2495 = _T_75183 ? _T_35064 : _GEN_345;
  assign _T_75223 = _T_99474 & _T_35090;
  assign _GEN_2496 = _T_75223 ? _T_35104 : _GEN_346;
  assign _T_75263 = _T_99474 & _T_35130;
  assign _GEN_2497 = _T_75263 ? _T_35144 : _GEN_347;
  assign _T_75303 = _T_99474 & _T_35170;
  assign _GEN_2498 = _T_75303 ? _T_35184 : _GEN_348;
  assign _GEN_7141 = {{8'd0}, _T_23996};
  assign _T_75399 = _GEN_7141 << 8;
  assign _GEN_7142 = {{8'd0}, _T_23994};
  assign _T_75403 = _GEN_7142 | _T_75399;
  assign _GEN_7143 = {{16'd0}, _T_23998};
  assign _T_75439 = _GEN_7143 << 16;
  assign _GEN_7144 = {{8'd0}, _T_75403};
  assign _T_75443 = _GEN_7144 | _T_75439;
  assign _GEN_7145 = {{24'd0}, _T_24000};
  assign _T_75479 = _GEN_7145 << 24;
  assign _GEN_7146 = {{8'd0}, _T_75443};
  assign _T_75483 = _GEN_7146 | _T_75479;
  assign _GEN_7147 = {{8'd0}, _T_24100};
  assign _T_75559 = _GEN_7147 << 8;
  assign _GEN_7148 = {{8'd0}, _T_24098};
  assign _T_75563 = _GEN_7148 | _T_75559;
  assign _GEN_7149 = {{16'd0}, _T_24102};
  assign _T_75599 = _GEN_7149 << 16;
  assign _GEN_7150 = {{8'd0}, _T_75563};
  assign _T_75603 = _GEN_7150 | _T_75599;
  assign _GEN_7151 = {{24'd0}, _T_24104};
  assign _T_75639 = _GEN_7151 << 24;
  assign _GEN_7152 = {{8'd0}, _T_75603};
  assign _T_75643 = _GEN_7152 | _T_75639;
  assign _GEN_7153 = {{8'd0}, _T_25276};
  assign _T_75719 = _GEN_7153 << 8;
  assign _GEN_7154 = {{8'd0}, _T_25274};
  assign _T_75723 = _GEN_7154 | _T_75719;
  assign _GEN_7155 = {{16'd0}, _T_25278};
  assign _T_75759 = _GEN_7155 << 16;
  assign _GEN_7156 = {{8'd0}, _T_75723};
  assign _T_75763 = _GEN_7156 | _T_75759;
  assign _GEN_7157 = {{24'd0}, _T_25280};
  assign _T_75799 = _GEN_7157 << 24;
  assign _GEN_7158 = {{8'd0}, _T_75763};
  assign _T_75803 = _GEN_7158 | _T_75799;
  assign _GEN_7159 = {{8'd0}, _T_24220};
  assign _T_75879 = _GEN_7159 << 8;
  assign _GEN_7160 = {{8'd0}, _T_24218};
  assign _T_75883 = _GEN_7160 | _T_75879;
  assign _GEN_7161 = {{16'd0}, _T_24222};
  assign _T_75919 = _GEN_7161 << 16;
  assign _GEN_7162 = {{8'd0}, _T_75883};
  assign _T_75923 = _GEN_7162 | _T_75919;
  assign _GEN_7163 = {{24'd0}, _T_24224};
  assign _T_75959 = _GEN_7163 << 24;
  assign _GEN_7164 = {{8'd0}, _T_75923};
  assign _T_75963 = _GEN_7164 | _T_75959;
  assign _GEN_7165 = {{8'd0}, _T_25156};
  assign _T_76039 = _GEN_7165 << 8;
  assign _GEN_7166 = {{8'd0}, _T_25154};
  assign _T_76043 = _GEN_7166 | _T_76039;
  assign _GEN_7167 = {{16'd0}, _T_25158};
  assign _T_76079 = _GEN_7167 << 16;
  assign _GEN_7168 = {{8'd0}, _T_76043};
  assign _T_76083 = _GEN_7168 | _T_76079;
  assign _GEN_7169 = {{24'd0}, _T_25160};
  assign _T_76119 = _GEN_7169 << 24;
  assign _GEN_7170 = {{8'd0}, _T_76083};
  assign _T_76123 = _GEN_7170 | _T_76119;
  assign _GEN_7171 = {{8'd0}, _T_24980};
  assign _T_76199 = _GEN_7171 << 8;
  assign _GEN_7172 = {{8'd0}, _T_24978};
  assign _T_76203 = _GEN_7172 | _T_76199;
  assign _GEN_7173 = {{16'd0}, _T_24982};
  assign _T_76239 = _GEN_7173 << 16;
  assign _GEN_7174 = {{8'd0}, _T_76203};
  assign _T_76243 = _GEN_7174 | _T_76239;
  assign _GEN_7175 = {{24'd0}, _T_24984};
  assign _T_76279 = _GEN_7175 << 24;
  assign _GEN_7176 = {{8'd0}, _T_76243};
  assign _T_76283 = _GEN_7176 | _T_76279;
  assign _GEN_7177 = {{8'd0}, _T_23796};
  assign _T_76359 = _GEN_7177 << 8;
  assign _GEN_7178 = {{8'd0}, _T_23794};
  assign _T_76363 = _GEN_7178 | _T_76359;
  assign _GEN_7179 = {{16'd0}, _T_23798};
  assign _T_76399 = _GEN_7179 << 16;
  assign _GEN_7180 = {{8'd0}, _T_76363};
  assign _T_76403 = _GEN_7180 | _T_76399;
  assign _GEN_7181 = {{24'd0}, _T_23800};
  assign _T_76439 = _GEN_7181 << 24;
  assign _GEN_7182 = {{8'd0}, _T_76403};
  assign _T_76443 = _GEN_7182 | _T_76439;
  assign _GEN_7183 = {{8'd0}, _T_24940};
  assign _T_76519 = _GEN_7183 << 8;
  assign _GEN_7184 = {{8'd0}, _T_24938};
  assign _T_76523 = _GEN_7184 | _T_76519;
  assign _GEN_7185 = {{16'd0}, _T_24942};
  assign _T_76559 = _GEN_7185 << 16;
  assign _GEN_7186 = {{8'd0}, _T_76523};
  assign _T_76563 = _GEN_7186 | _T_76559;
  assign _GEN_7187 = {{24'd0}, _T_24944};
  assign _T_76599 = _GEN_7187 << 24;
  assign _GEN_7188 = {{8'd0}, _T_76563};
  assign _T_76603 = _GEN_7188 | _T_76599;
  assign _GEN_7189 = {{8'd0}, _T_25076};
  assign _T_76679 = _GEN_7189 << 8;
  assign _GEN_7190 = {{8'd0}, _T_25074};
  assign _T_76683 = _GEN_7190 | _T_76679;
  assign _GEN_7191 = {{16'd0}, _T_25078};
  assign _T_76719 = _GEN_7191 << 16;
  assign _GEN_7192 = {{8'd0}, _T_76683};
  assign _T_76723 = _GEN_7192 | _T_76719;
  assign _GEN_7193 = {{24'd0}, _T_25080};
  assign _T_76759 = _GEN_7193 << 24;
  assign _GEN_7194 = {{8'd0}, _T_76723};
  assign _T_76763 = _GEN_7194 | _T_76759;
  assign _GEN_7195 = {{8'd0}, _T_23884};
  assign _T_76839 = _GEN_7195 << 8;
  assign _GEN_7196 = {{8'd0}, _T_23882};
  assign _T_76843 = _GEN_7196 | _T_76839;
  assign _GEN_7197 = {{16'd0}, _T_23886};
  assign _T_76879 = _GEN_7197 << 16;
  assign _GEN_7198 = {{8'd0}, _T_76843};
  assign _T_76883 = _GEN_7198 | _T_76879;
  assign _GEN_7199 = {{24'd0}, _T_23888};
  assign _T_76919 = _GEN_7199 << 24;
  assign _GEN_7200 = {{8'd0}, _T_76883};
  assign _T_76923 = _GEN_7200 | _T_76919;
  assign _GEN_7201 = {{8'd0}, _T_24684};
  assign _T_76999 = _GEN_7201 << 8;
  assign _GEN_7202 = {{8'd0}, _T_24682};
  assign _T_77003 = _GEN_7202 | _T_76999;
  assign _GEN_7203 = {{16'd0}, _T_24686};
  assign _T_77039 = _GEN_7203 << 16;
  assign _GEN_7204 = {{8'd0}, _T_77003};
  assign _T_77043 = _GEN_7204 | _T_77039;
  assign _GEN_7205 = {{24'd0}, _T_24688};
  assign _T_77079 = _GEN_7205 << 24;
  assign _GEN_7206 = {{8'd0}, _T_77043};
  assign _T_77083 = _GEN_7206 | _T_77079;
  assign _GEN_7207 = {{8'd0}, _T_24140};
  assign _T_77159 = _GEN_7207 << 8;
  assign _GEN_7208 = {{8'd0}, _T_24138};
  assign _T_77163 = _GEN_7208 | _T_77159;
  assign _GEN_7209 = {{16'd0}, _T_24142};
  assign _T_77199 = _GEN_7209 << 16;
  assign _GEN_7210 = {{8'd0}, _T_77163};
  assign _T_77203 = _GEN_7210 | _T_77199;
  assign _GEN_7211 = {{24'd0}, _T_24144};
  assign _T_77239 = _GEN_7211 << 24;
  assign _GEN_7212 = {{8'd0}, _T_77203};
  assign _T_77243 = _GEN_7212 | _T_77239;
  assign _T_77263 = _T_99442 & _T_35050;
  assign _GEN_2499 = _T_77263 ? _T_35064 : _GEN_329;
  assign _T_77303 = _T_99442 & _T_35090;
  assign _GEN_2500 = _T_77303 ? _T_35104 : _GEN_330;
  assign _T_77343 = _T_99442 & _T_35130;
  assign _GEN_2501 = _T_77343 ? _T_35144 : _GEN_331;
  assign _T_77383 = _T_99442 & _T_35170;
  assign _GEN_2502 = _T_77383 ? _T_35184 : _GEN_332;
  assign _GEN_7219 = {{8'd0}, _T_24308};
  assign _T_77479 = _GEN_7219 << 8;
  assign _GEN_7220 = {{8'd0}, _T_24306};
  assign _T_77483 = _GEN_7220 | _T_77479;
  assign _GEN_7221 = {{16'd0}, _T_24310};
  assign _T_77519 = _GEN_7221 << 16;
  assign _GEN_7222 = {{8'd0}, _T_77483};
  assign _T_77523 = _GEN_7222 | _T_77519;
  assign _GEN_7223 = {{24'd0}, _T_24312};
  assign _T_77559 = _GEN_7223 << 24;
  assign _GEN_7224 = {{8'd0}, _T_77523};
  assign _T_77563 = _GEN_7224 | _T_77559;
  assign _GEN_7225 = {{8'd0}, _T_24052};
  assign _T_77639 = _GEN_7225 << 8;
  assign _GEN_7226 = {{8'd0}, _T_24050};
  assign _T_77643 = _GEN_7226 | _T_77639;
  assign _GEN_7227 = {{16'd0}, _T_24054};
  assign _T_77679 = _GEN_7227 << 16;
  assign _GEN_7228 = {{8'd0}, _T_77643};
  assign _T_77683 = _GEN_7228 | _T_77679;
  assign _GEN_7229 = {{24'd0}, _T_24056};
  assign _T_77719 = _GEN_7229 << 24;
  assign _GEN_7230 = {{8'd0}, _T_77683};
  assign _T_77723 = _GEN_7230 | _T_77719;
  assign _GEN_7231 = {{8'd0}, _T_24428};
  assign _T_77799 = _GEN_7231 << 8;
  assign _GEN_7232 = {{8'd0}, _T_24426};
  assign _T_77803 = _GEN_7232 | _T_77799;
  assign _GEN_7233 = {{16'd0}, _T_24430};
  assign _T_77839 = _GEN_7233 << 16;
  assign _GEN_7234 = {{8'd0}, _T_77803};
  assign _T_77843 = _GEN_7234 | _T_77839;
  assign _GEN_7235 = {{24'd0}, _T_24432};
  assign _T_77879 = _GEN_7235 << 24;
  assign _GEN_7236 = {{8'd0}, _T_77843};
  assign _T_77883 = _GEN_7236 | _T_77879;
  assign _GEN_7237 = {{8'd0}, _T_25748};
  assign _T_77959 = _GEN_7237 << 8;
  assign _GEN_7238 = {{8'd0}, _T_25746};
  assign _T_77963 = _GEN_7238 | _T_77959;
  assign _GEN_7239 = {{16'd0}, _T_25750};
  assign _T_77999 = _GEN_7239 << 16;
  assign _GEN_7240 = {{8'd0}, _T_77963};
  assign _T_78003 = _GEN_7240 | _T_77999;
  assign _GEN_7241 = {{24'd0}, _T_25752};
  assign _T_78039 = _GEN_7241 << 24;
  assign _GEN_7242 = {{8'd0}, _T_78003};
  assign _T_78043 = _GEN_7242 | _T_78039;
  assign _GEN_7243 = {{8'd0}, _T_23844};
  assign _T_78119 = _GEN_7243 << 8;
  assign _GEN_7244 = {{8'd0}, _T_23842};
  assign _T_78123 = _GEN_7244 | _T_78119;
  assign _GEN_7245 = {{16'd0}, _T_23846};
  assign _T_78159 = _GEN_7245 << 16;
  assign _GEN_7246 = {{8'd0}, _T_78123};
  assign _T_78163 = _GEN_7246 | _T_78159;
  assign _GEN_7247 = {{24'd0}, _T_23848};
  assign _T_78199 = _GEN_7247 << 24;
  assign _GEN_7248 = {{8'd0}, _T_78163};
  assign _T_78203 = _GEN_7248 | _T_78199;
  assign _GEN_7249 = {{8'd0}, _T_24564};
  assign _T_78279 = _GEN_7249 << 8;
  assign _GEN_7250 = {{8'd0}, _T_24562};
  assign _T_78283 = _GEN_7250 | _T_78279;
  assign _GEN_7251 = {{16'd0}, _T_24566};
  assign _T_78319 = _GEN_7251 << 16;
  assign _GEN_7252 = {{8'd0}, _T_78283};
  assign _T_78323 = _GEN_7252 | _T_78319;
  assign _GEN_7253 = {{24'd0}, _T_24568};
  assign _T_78359 = _GEN_7253 << 24;
  assign _GEN_7254 = {{8'd0}, _T_78323};
  assign _T_78363 = _GEN_7254 | _T_78359;
  assign _GEN_7255 = {{8'd0}, _T_25196};
  assign _T_78439 = _GEN_7255 << 8;
  assign _GEN_7256 = {{8'd0}, _T_25194};
  assign _T_78443 = _GEN_7256 | _T_78439;
  assign _GEN_7257 = {{16'd0}, _T_25198};
  assign _T_78479 = _GEN_7257 << 16;
  assign _GEN_7258 = {{8'd0}, _T_78443};
  assign _T_78483 = _GEN_7258 | _T_78479;
  assign _GEN_7259 = {{24'd0}, _T_25200};
  assign _T_78519 = _GEN_7259 << 24;
  assign _GEN_7260 = {{8'd0}, _T_78483};
  assign _T_78523 = _GEN_7260 | _T_78519;
  assign _GEN_7261 = {{8'd0}, _T_25492};
  assign _T_78599 = _GEN_7261 << 8;
  assign _GEN_7262 = {{8'd0}, _T_25490};
  assign _T_78603 = _GEN_7262 | _T_78599;
  assign _GEN_7263 = {{16'd0}, _T_25494};
  assign _T_78639 = _GEN_7263 << 16;
  assign _GEN_7264 = {{8'd0}, _T_78603};
  assign _T_78643 = _GEN_7264 | _T_78639;
  assign _GEN_7265 = {{24'd0}, _T_25496};
  assign _T_78679 = _GEN_7265 << 24;
  assign _GEN_7266 = {{8'd0}, _T_78643};
  assign _T_78683 = _GEN_7266 | _T_78679;
  assign _GEN_7267 = {{8'd0}, _T_24900};
  assign _T_78759 = _GEN_7267 << 8;
  assign _GEN_7268 = {{8'd0}, _T_24898};
  assign _T_78763 = _GEN_7268 | _T_78759;
  assign _GEN_7269 = {{16'd0}, _T_24902};
  assign _T_78799 = _GEN_7269 << 16;
  assign _GEN_7270 = {{8'd0}, _T_78763};
  assign _T_78803 = _GEN_7270 | _T_78799;
  assign _GEN_7271 = {{24'd0}, _T_24904};
  assign _T_78839 = _GEN_7271 << 24;
  assign _GEN_7272 = {{8'd0}, _T_78803};
  assign _T_78843 = _GEN_7272 | _T_78839;
  assign _GEN_7273 = {{8'd0}, _T_23964};
  assign _T_79079 = _GEN_7273 << 8;
  assign _GEN_7274 = {{8'd0}, _T_23962};
  assign _T_79083 = _GEN_7274 | _T_79079;
  assign _GEN_7275 = {{16'd0}, _T_23966};
  assign _T_79119 = _GEN_7275 << 16;
  assign _GEN_7276 = {{8'd0}, _T_79083};
  assign _T_79123 = _GEN_7276 | _T_79119;
  assign _GEN_7277 = {{24'd0}, _T_23968};
  assign _T_79159 = _GEN_7277 << 24;
  assign _GEN_7278 = {{8'd0}, _T_79123};
  assign _T_79163 = _GEN_7278 | _T_79159;
  assign _GEN_7279 = {{8'd0}, _T_25020};
  assign _T_79239 = _GEN_7279 << 8;
  assign _GEN_7280 = {{8'd0}, _T_25018};
  assign _T_79243 = _GEN_7280 | _T_79239;
  assign _GEN_7281 = {{16'd0}, _T_25022};
  assign _T_79279 = _GEN_7281 << 16;
  assign _GEN_7282 = {{8'd0}, _T_79243};
  assign _T_79283 = _GEN_7282 | _T_79279;
  assign _GEN_7283 = {{24'd0}, _T_25024};
  assign _T_79319 = _GEN_7283 << 24;
  assign _GEN_7284 = {{8'd0}, _T_79283};
  assign _T_79323 = _GEN_7284 | _T_79319;
  assign _GEN_7285 = {{8'd0}, _T_24860};
  assign _T_79399 = _GEN_7285 << 8;
  assign _GEN_7286 = {{8'd0}, _T_24858};
  assign _T_79403 = _GEN_7286 | _T_79399;
  assign _GEN_7287 = {{16'd0}, _T_24862};
  assign _T_79439 = _GEN_7287 << 16;
  assign _GEN_7288 = {{8'd0}, _T_79403};
  assign _T_79443 = _GEN_7288 | _T_79439;
  assign _GEN_7289 = {{24'd0}, _T_24864};
  assign _T_79479 = _GEN_7289 << 24;
  assign _GEN_7290 = {{8'd0}, _T_79443};
  assign _T_79483 = _GEN_7290 | _T_79479;
  assign _GEN_7291 = {{8'd0}, _T_25412};
  assign _T_79559 = _GEN_7291 << 8;
  assign _GEN_7292 = {{8'd0}, _T_25410};
  assign _T_79563 = _GEN_7292 | _T_79559;
  assign _GEN_7293 = {{16'd0}, _T_25414};
  assign _T_79599 = _GEN_7293 << 16;
  assign _GEN_7294 = {{8'd0}, _T_79563};
  assign _T_79603 = _GEN_7294 | _T_79599;
  assign _GEN_7295 = {{24'd0}, _T_25416};
  assign _T_79639 = _GEN_7295 << 24;
  assign _GEN_7296 = {{8'd0}, _T_79603};
  assign _T_79643 = _GEN_7296 | _T_79639;
  assign _GEN_7297 = {{8'd0}, _T_24356};
  assign _T_79719 = _GEN_7297 << 8;
  assign _GEN_7298 = {{8'd0}, _T_24354};
  assign _T_79723 = _GEN_7298 | _T_79719;
  assign _GEN_7299 = {{16'd0}, _T_24358};
  assign _T_79759 = _GEN_7299 << 16;
  assign _GEN_7300 = {{8'd0}, _T_79723};
  assign _T_79763 = _GEN_7300 | _T_79759;
  assign _GEN_7301 = {{24'd0}, _T_24360};
  assign _T_79799 = _GEN_7301 << 24;
  assign _GEN_7302 = {{8'd0}, _T_79763};
  assign _T_79803 = _GEN_7302 | _T_79799;
  assign _GEN_7303 = {{8'd0}, _T_25116};
  assign _T_79879 = _GEN_7303 << 8;
  assign _GEN_7304 = {{8'd0}, _T_25114};
  assign _T_79883 = _GEN_7304 | _T_79879;
  assign _GEN_7305 = {{16'd0}, _T_25118};
  assign _T_79919 = _GEN_7305 << 16;
  assign _GEN_7306 = {{8'd0}, _T_79883};
  assign _T_79923 = _GEN_7306 | _T_79919;
  assign _GEN_7307 = {{24'd0}, _T_25120};
  assign _T_79959 = _GEN_7307 << 24;
  assign _GEN_7308 = {{8'd0}, _T_79923};
  assign _T_79963 = _GEN_7308 | _T_79959;
  assign _GEN_7309 = {{8'd0}, _T_25372};
  assign _T_80199 = _GEN_7309 << 8;
  assign _GEN_7310 = {{8'd0}, _T_25370};
  assign _T_80203 = _GEN_7310 | _T_80199;
  assign _GEN_7311 = {{16'd0}, _T_25374};
  assign _T_80239 = _GEN_7311 << 16;
  assign _GEN_7312 = {{8'd0}, _T_80203};
  assign _T_80243 = _GEN_7312 | _T_80239;
  assign _GEN_7313 = {{24'd0}, _T_25376};
  assign _T_80279 = _GEN_7313 << 24;
  assign _GEN_7314 = {{8'd0}, _T_80243};
  assign _T_80283 = _GEN_7314 | _T_80279;
  assign _GEN_7315 = {{8'd0}, _T_23916};
  assign _T_80359 = _GEN_7315 << 8;
  assign _GEN_7316 = {{8'd0}, _T_23914};
  assign _T_80363 = _GEN_7316 | _T_80359;
  assign _GEN_7317 = {{16'd0}, _T_23918};
  assign _T_80399 = _GEN_7317 << 16;
  assign _GEN_7318 = {{8'd0}, _T_80363};
  assign _T_80403 = _GEN_7318 | _T_80399;
  assign _GEN_7319 = {{24'd0}, _T_23920};
  assign _T_80439 = _GEN_7319 << 24;
  assign _GEN_7320 = {{8'd0}, _T_80403};
  assign _T_80443 = _GEN_7320 | _T_80439;
  assign _GEN_7321 = {{8'd0}, _T_25236};
  assign _T_80519 = _GEN_7321 << 8;
  assign _GEN_7322 = {{8'd0}, _T_25234};
  assign _T_80523 = _GEN_7322 | _T_80519;
  assign _GEN_7323 = {{16'd0}, _T_25238};
  assign _T_80559 = _GEN_7323 << 16;
  assign _GEN_7324 = {{8'd0}, _T_80523};
  assign _T_80563 = _GEN_7324 | _T_80559;
  assign _GEN_7325 = {{24'd0}, _T_25240};
  assign _T_80599 = _GEN_7325 << 24;
  assign _GEN_7326 = {{8'd0}, _T_80563};
  assign _T_80603 = _GEN_7326 | _T_80599;
  assign _GEN_7327 = {{8'd0}, _T_25708};
  assign _T_80679 = _GEN_7327 << 8;
  assign _GEN_7328 = {{8'd0}, _T_25706};
  assign _T_80683 = _GEN_7328 | _T_80679;
  assign _GEN_7329 = {{16'd0}, _T_25710};
  assign _T_80719 = _GEN_7329 << 16;
  assign _GEN_7330 = {{8'd0}, _T_80683};
  assign _T_80723 = _GEN_7330 | _T_80719;
  assign _GEN_7331 = {{24'd0}, _T_25712};
  assign _T_80759 = _GEN_7331 << 24;
  assign _GEN_7332 = {{8'd0}, _T_80723};
  assign _T_80763 = _GEN_7332 | _T_80759;
  assign _GEN_7333 = {{8'd0}, _T_24652};
  assign _T_80839 = _GEN_7333 << 8;
  assign _GEN_7334 = {{8'd0}, _T_24650};
  assign _T_80843 = _GEN_7334 | _T_80839;
  assign _GEN_7335 = {{16'd0}, _T_24654};
  assign _T_80879 = _GEN_7335 << 16;
  assign _GEN_7336 = {{8'd0}, _T_80843};
  assign _T_80883 = _GEN_7336 | _T_80879;
  assign _GEN_7337 = {{24'd0}, _T_24656};
  assign _T_80919 = _GEN_7337 << 24;
  assign _GEN_7338 = {{8'd0}, _T_80883};
  assign _T_80923 = _GEN_7338 | _T_80919;
  assign _GEN_7339 = {{8'd0}, _T_24276};
  assign _T_80999 = _GEN_7339 << 8;
  assign _GEN_7340 = {{8'd0}, _T_24274};
  assign _T_81003 = _GEN_7340 | _T_80999;
  assign _GEN_7341 = {{16'd0}, _T_24278};
  assign _T_81039 = _GEN_7341 << 16;
  assign _GEN_7342 = {{8'd0}, _T_81003};
  assign _T_81043 = _GEN_7342 | _T_81039;
  assign _GEN_7343 = {{24'd0}, _T_24280};
  assign _T_81079 = _GEN_7343 << 24;
  assign _GEN_7344 = {{8'd0}, _T_81043};
  assign _T_81083 = _GEN_7344 | _T_81079;
  assign _GEN_7345 = {{8'd0}, _T_25588};
  assign _T_81159 = _GEN_7345 << 8;
  assign _GEN_7346 = {{8'd0}, _T_25586};
  assign _T_81163 = _GEN_7346 | _T_81159;
  assign _GEN_7347 = {{16'd0}, _T_25590};
  assign _T_81199 = _GEN_7347 << 16;
  assign _GEN_7348 = {{8'd0}, _T_81163};
  assign _T_81203 = _GEN_7348 | _T_81199;
  assign _GEN_7349 = {{24'd0}, _T_25592};
  assign _T_81239 = _GEN_7349 << 24;
  assign _GEN_7350 = {{8'd0}, _T_81203};
  assign _T_81243 = _GEN_7350 | _T_81239;
  assign _GEN_7351 = {{8'd0}, _T_24396};
  assign _T_81319 = _GEN_7351 << 8;
  assign _GEN_7352 = {{8'd0}, _T_24394};
  assign _T_81323 = _GEN_7352 | _T_81319;
  assign _GEN_7353 = {{16'd0}, _T_24398};
  assign _T_81359 = _GEN_7353 << 16;
  assign _GEN_7354 = {{8'd0}, _T_81323};
  assign _T_81363 = _GEN_7354 | _T_81359;
  assign _GEN_7355 = {{24'd0}, _T_24400};
  assign _T_81399 = _GEN_7355 << 24;
  assign _GEN_7356 = {{8'd0}, _T_81363};
  assign _T_81403 = _GEN_7356 | _T_81399;
  assign _GEN_7357 = {{8'd0}, _T_25452};
  assign _T_81479 = _GEN_7357 << 8;
  assign _GEN_7358 = {{8'd0}, _T_25450};
  assign _T_81483 = _GEN_7358 | _T_81479;
  assign _GEN_7359 = {{16'd0}, _T_25454};
  assign _T_81519 = _GEN_7359 << 16;
  assign _GEN_7360 = {{8'd0}, _T_81483};
  assign _T_81523 = _GEN_7360 | _T_81519;
  assign _GEN_7361 = {{24'd0}, _T_25456};
  assign _T_81559 = _GEN_7361 << 24;
  assign _GEN_7362 = {{8'd0}, _T_81523};
  assign _T_81563 = _GEN_7362 | _T_81559;
  assign _GEN_7363 = {{8'd0}, _T_24532};
  assign _T_81639 = _GEN_7363 << 8;
  assign _GEN_7364 = {{8'd0}, _T_24530};
  assign _T_81643 = _GEN_7364 | _T_81639;
  assign _GEN_7365 = {{16'd0}, _T_24534};
  assign _T_81679 = _GEN_7365 << 16;
  assign _GEN_7366 = {{8'd0}, _T_81643};
  assign _T_81683 = _GEN_7366 | _T_81679;
  assign _GEN_7367 = {{24'd0}, _T_24536};
  assign _T_81719 = _GEN_7367 << 24;
  assign _GEN_7368 = {{8'd0}, _T_81683};
  assign _T_81723 = _GEN_7368 | _T_81719;
  assign _GEN_7369 = {{8'd0}, _T_24172};
  assign _T_81799 = _GEN_7369 << 8;
  assign _GEN_7370 = {{8'd0}, _T_24170};
  assign _T_81803 = _GEN_7370 | _T_81799;
  assign _GEN_7371 = {{16'd0}, _T_24174};
  assign _T_81839 = _GEN_7371 << 16;
  assign _GEN_7372 = {{8'd0}, _T_81803};
  assign _T_81843 = _GEN_7372 | _T_81839;
  assign _GEN_7373 = {{24'd0}, _T_24176};
  assign _T_81879 = _GEN_7373 << 24;
  assign _GEN_7374 = {{8'd0}, _T_81843};
  assign _T_81883 = _GEN_7374 | _T_81879;
  assign _T_81903 = _T_99482 & _T_35050;
  assign _GEN_2503 = _T_81903 ? _T_35064 : _GEN_349;
  assign _T_81943 = _T_99482 & _T_35090;
  assign _GEN_2504 = _T_81943 ? _T_35104 : _GEN_350;
  assign _T_81983 = _T_99482 & _T_35130;
  assign _GEN_2505 = _T_81983 ? _T_35144 : _GEN_351;
  assign _T_82023 = _T_99482 & _T_35170;
  assign _GEN_2506 = _T_82023 ? _T_35184 : _GEN_352;
  assign _GEN_7381 = {{8'd0}, _T_25628};
  assign _T_82119 = _GEN_7381 << 8;
  assign _GEN_7382 = {{8'd0}, _T_25626};
  assign _T_82123 = _GEN_7382 | _T_82119;
  assign _GEN_7383 = {{16'd0}, _T_25630};
  assign _T_82159 = _GEN_7383 << 16;
  assign _GEN_7384 = {{8'd0}, _T_82123};
  assign _T_82163 = _GEN_7384 | _T_82159;
  assign _GEN_7385 = {{24'd0}, _T_25632};
  assign _T_82199 = _GEN_7385 << 24;
  assign _GEN_7386 = {{8'd0}, _T_82163};
  assign _T_82203 = _GEN_7386 | _T_82199;
  assign _T_82223 = _T_99538 & _T_35050;
  assign _GEN_2507 = _T_82223 ? _T_35064 : _GEN_377;
  assign _T_82263 = _T_99538 & _T_35090;
  assign _GEN_2508 = _T_82263 ? _T_35104 : _GEN_378;
  assign _T_82303 = _T_99538 & _T_35130;
  assign _GEN_2509 = _T_82303 ? _T_35144 : _GEN_379;
  assign _T_82343 = _T_99538 & _T_35170;
  assign _GEN_2510 = _T_82343 ? _T_35184 : _GEN_380;
  assign _GEN_7393 = {{8'd0}, _T_25668};
  assign _T_82439 = _GEN_7393 << 8;
  assign _GEN_7394 = {{8'd0}, _T_25666};
  assign _T_82443 = _GEN_7394 | _T_82439;
  assign _GEN_7395 = {{16'd0}, _T_25670};
  assign _T_82479 = _GEN_7395 << 16;
  assign _GEN_7396 = {{8'd0}, _T_82443};
  assign _T_82483 = _GEN_7396 | _T_82479;
  assign _GEN_7397 = {{24'd0}, _T_25672};
  assign _T_82519 = _GEN_7397 << 24;
  assign _GEN_7398 = {{8'd0}, _T_82483};
  assign _T_82523 = _GEN_7398 | _T_82519;
  assign _GEN_7399 = {{8'd0}, _T_25332};
  assign _T_82599 = _GEN_7399 << 8;
  assign _GEN_7400 = {{8'd0}, _T_25330};
  assign _T_82603 = _GEN_7400 | _T_82599;
  assign _GEN_7401 = {{16'd0}, _T_25334};
  assign _T_82639 = _GEN_7401 << 16;
  assign _GEN_7402 = {{8'd0}, _T_82603};
  assign _T_82643 = _GEN_7402 | _T_82639;
  assign _GEN_7403 = {{24'd0}, _T_25336};
  assign _T_82679 = _GEN_7403 << 24;
  assign _GEN_7404 = {{8'd0}, _T_82643};
  assign _T_82683 = _GEN_7404 | _T_82679;
  assign _GEN_7405 = {{8'd0}, _T_24612};
  assign _T_82759 = _GEN_7405 << 8;
  assign _GEN_7406 = {{8'd0}, _T_24610};
  assign _T_82763 = _GEN_7406 | _T_82759;
  assign _GEN_7407 = {{16'd0}, _T_24614};
  assign _T_82799 = _GEN_7407 << 16;
  assign _GEN_7408 = {{8'd0}, _T_82763};
  assign _T_82803 = _GEN_7408 | _T_82799;
  assign _GEN_7409 = {{24'd0}, _T_24616};
  assign _T_82839 = _GEN_7409 << 24;
  assign _GEN_7410 = {{8'd0}, _T_82803};
  assign _T_82843 = _GEN_7410 | _T_82839;
  assign _T_82844 = _T_25900[0];
  assign _T_82845 = _T_25900[1];
  assign _T_82846 = _T_25900[2];
  assign _T_82847 = _T_25900[3];
  assign _T_82848 = _T_25900[4];
  assign _T_82849 = _T_25900[5];
  assign _T_82850 = _T_25900[6];
  assign _T_82851 = _T_25900[7];
  assign _T_82852 = _T_25900[8];
  assign _T_82854 = {_T_82845,_T_82844};
  assign _T_82855 = {_T_82847,_T_82846};
  assign _T_82856 = {_T_82855,_T_82854};
  assign _T_82857 = {_T_82849,_T_82848};
  assign _T_82858 = {_T_82852,_T_82851};
  assign _T_82859 = {_T_82858,_T_82850};
  assign _T_82860 = {_T_82859,_T_82857};
  assign _T_82861 = {_T_82860,_T_82856};
  assign _T_82881 = 512'h1 << _T_82861;
  assign _T_82946 = _T_82881[64];
  assign _T_82947 = _T_82881[65];
  assign _T_82948 = _T_82881[66];
  assign _T_82949 = _T_82881[67];
  assign _T_83090 = _T_82881[208];
  assign _T_83091 = _T_82881[209];
  assign _T_83092 = _T_82881[210];
  assign _T_83093 = _T_82881[211];
  assign _T_83094 = _T_82881[212];
  assign _T_83095 = _T_82881[213];
  assign _T_83096 = _T_82881[214];
  assign _T_83097 = _T_82881[215];
  assign _T_83098 = _T_82881[216];
  assign _T_83099 = _T_82881[217];
  assign _T_83100 = _T_82881[218];
  assign _T_83101 = _T_82881[219];
  assign _T_83102 = _T_82881[220];
  assign _T_83103 = _T_82881[221];
  assign _T_83104 = _T_82881[222];
  assign _T_83105 = _T_82881[223];
  assign _T_83106 = _T_82881[224];
  assign _T_83908 = io_hart_in_0_a_valid & io_hart_in_0_d_ready;
  assign _T_88525 = _T_25899 == 1'h0;
  assign _T_88526 = _T_83908 & _T_88525;
  assign _T_89041 = _T_88526 & _T_82946;
  assign _T_89049 = _T_88526 & _T_82947;
  assign _T_89057 = _T_88526 & _T_82948;
  assign _T_89065 = _T_88526 & _T_82949;
  assign _T_90193 = _T_88526 & _T_83090;
  assign _T_90201 = _T_88526 & _T_83091;
  assign _T_90209 = _T_88526 & _T_83092;
  assign _T_90217 = _T_88526 & _T_83093;
  assign _T_90225 = _T_88526 & _T_83094;
  assign _T_90233 = _T_88526 & _T_83095;
  assign _T_90241 = _T_88526 & _T_83096;
  assign _T_90249 = _T_88526 & _T_83097;
  assign _T_90257 = _T_88526 & _T_83098;
  assign _T_90265 = _T_88526 & _T_83099;
  assign _T_90273 = _T_88526 & _T_83100;
  assign _T_90281 = _T_88526 & _T_83101;
  assign _T_90289 = _T_88526 & _T_83102;
  assign _T_90297 = _T_88526 & _T_83103;
  assign _T_90305 = _T_88526 & _T_83104;
  assign _T_90313 = _T_88526 & _T_83105;
  assign _T_90321 = _T_88526 & _T_83106;
  assign _T_98274 = _T_89041 & _T_28219;
  assign _T_98282 = _T_89049 & _T_27814;
  assign _T_98290 = _T_89057 & _T_28597;
  assign _T_98298 = _T_89065 & _T_28903;
  assign _T_99426 = _T_90193 & _T_28498;
  assign _T_99434 = _T_90201 & _T_28777;
  assign _T_99442 = _T_90209 & _T_29371;
  assign _T_99450 = _T_90217 & _T_27409;
  assign _T_99458 = _T_90225 & _T_28039;
  assign _T_99466 = _T_90233 & _T_28570;
  assign _T_99474 = _T_90241 & _T_29254;
  assign _T_99482 = _T_90249 & _T_29632;
  assign _T_99490 = _T_90257 & _T_27355;
  assign _T_99498 = _T_90265 & _T_27040;
  assign _T_99506 = _T_90273 & _T_29083;
  assign _T_99514 = _T_90281 & _T_28399;
  assign _T_99522 = _T_90289 & _T_27661;
  assign _T_99530 = _T_90297 & _T_27481;
  assign _T_99538 = _T_90305 & _T_29650;
  assign _T_99546 = _T_90313 & _T_28660;
  assign _T_99554 = _T_90321 & _T_27895;
  assign _T_102902_64 = {{22'd0}, _T_50184};
  assign _T_102902_65 = {{22'd0}, _T_50184};
  assign _T_102902_66 = {{22'd0}, _T_50184};
  assign _T_102902_67 = {{22'd0}, _T_50184};
  assign _GEN_4555 = 9'h1 == _T_82861 ? _T_28183 : _T_27616;
  assign _GEN_4556 = 9'h2 == _T_82861 ? _T_27427 : _GEN_4555;
  assign _GEN_4557 = 9'h3 == _T_82861 ? _T_28057 : _GEN_4556;
  assign _GEN_4558 = 9'h4 == _T_82861 ? _T_28795 : _GEN_4557;
  assign _GEN_4559 = 9'h5 == _T_82861 ? _T_29101 : _GEN_4558;
  assign _GEN_4560 = 9'h6 == _T_82861 ? _T_26986 : _GEN_4559;
  assign _GEN_4561 = 9'h7 == _T_82861 ? _T_27904 : _GEN_4560;
  assign _GEN_4562 = 9'h8 == _T_82861 ? _T_28588 : _GEN_4561;
  assign _GEN_4563 = 9'h9 == _T_82861 ? _T_28624 : _GEN_4562;
  assign _GEN_4564 = 9'ha == _T_82861 ? _T_27841 : _GEN_4563;
  assign _GEN_4565 = 9'hb == _T_82861 ? _T_27031 : _GEN_4564;
  assign _GEN_4566 = 9'hc == _T_82861 ? _T_29065 : _GEN_4565;
  assign _GEN_4567 = 9'hd == _T_82861 ? _T_28831 : _GEN_4566;
  assign _GEN_4568 = 9'he == _T_82861 ? _T_28021 : _GEN_4567;
  assign _GEN_4569 = 9'hf == _T_82861 ? _T_27553 : _GEN_4568;
  assign _GEN_4570 = 9'h10 == _T_82861 ? _T_29524 : _GEN_4569;
  assign _GEN_4571 = 9'h11 == _T_82861 ? _T_27643 : _GEN_4570;
  assign _GEN_4572 = 9'h12 == _T_82861 ? _T_28147 : _GEN_4571;
  assign _GEN_4573 = 9'h13 == _T_82861 ? _T_28759 : _GEN_4572;
  assign _GEN_4574 = 9'h14 == _T_82861 ? _T_29461 : _GEN_4573;
  assign _GEN_4575 = 9'h15 == _T_82861 ? _T_27130 : _GEN_4574;
  assign _GEN_4576 = 9'h16 == _T_82861 ? _T_27679 : _GEN_4575;
  assign _GEN_4577 = 9'h17 == _T_82861 ? _T_28552 : _GEN_4576;
  assign _GEN_4578 = 9'h18 == _T_82861 ? 1'h1 : _GEN_4577;
  assign _GEN_4579 = 9'h19 == _T_82861 ? 1'h1 : _GEN_4578;
  assign _GEN_4580 = 9'h1a == _T_82861 ? 1'h1 : _GEN_4579;
  assign _GEN_4581 = 9'h1b == _T_82861 ? 1'h1 : _GEN_4580;
  assign _GEN_4582 = 9'h1c == _T_82861 ? 1'h1 : _GEN_4581;
  assign _GEN_4583 = 9'h1d == _T_82861 ? 1'h1 : _GEN_4582;
  assign _GEN_4584 = 9'h1e == _T_82861 ? 1'h1 : _GEN_4583;
  assign _GEN_4585 = 9'h1f == _T_82861 ? 1'h1 : _GEN_4584;
  assign _GEN_4586 = 9'h20 == _T_82861 ? 1'h1 : _GEN_4585;
  assign _GEN_4587 = 9'h21 == _T_82861 ? 1'h1 : _GEN_4586;
  assign _GEN_4588 = 9'h22 == _T_82861 ? 1'h1 : _GEN_4587;
  assign _GEN_4589 = 9'h23 == _T_82861 ? 1'h1 : _GEN_4588;
  assign _GEN_4590 = 9'h24 == _T_82861 ? 1'h1 : _GEN_4589;
  assign _GEN_4591 = 9'h25 == _T_82861 ? 1'h1 : _GEN_4590;
  assign _GEN_4592 = 9'h26 == _T_82861 ? 1'h1 : _GEN_4591;
  assign _GEN_4593 = 9'h27 == _T_82861 ? 1'h1 : _GEN_4592;
  assign _GEN_4594 = 9'h28 == _T_82861 ? 1'h1 : _GEN_4593;
  assign _GEN_4595 = 9'h29 == _T_82861 ? 1'h1 : _GEN_4594;
  assign _GEN_4596 = 9'h2a == _T_82861 ? 1'h1 : _GEN_4595;
  assign _GEN_4597 = 9'h2b == _T_82861 ? 1'h1 : _GEN_4596;
  assign _GEN_4598 = 9'h2c == _T_82861 ? 1'h1 : _GEN_4597;
  assign _GEN_4599 = 9'h2d == _T_82861 ? 1'h1 : _GEN_4598;
  assign _GEN_4600 = 9'h2e == _T_82861 ? 1'h1 : _GEN_4599;
  assign _GEN_4601 = 9'h2f == _T_82861 ? 1'h1 : _GEN_4600;
  assign _GEN_4602 = 9'h30 == _T_82861 ? 1'h1 : _GEN_4601;
  assign _GEN_4603 = 9'h31 == _T_82861 ? 1'h1 : _GEN_4602;
  assign _GEN_4604 = 9'h32 == _T_82861 ? 1'h1 : _GEN_4603;
  assign _GEN_4605 = 9'h33 == _T_82861 ? 1'h1 : _GEN_4604;
  assign _GEN_4606 = 9'h34 == _T_82861 ? 1'h1 : _GEN_4605;
  assign _GEN_4607 = 9'h35 == _T_82861 ? 1'h1 : _GEN_4606;
  assign _GEN_4608 = 9'h36 == _T_82861 ? 1'h1 : _GEN_4607;
  assign _GEN_4609 = 9'h37 == _T_82861 ? 1'h1 : _GEN_4608;
  assign _GEN_4610 = 9'h38 == _T_82861 ? 1'h1 : _GEN_4609;
  assign _GEN_4611 = 9'h39 == _T_82861 ? 1'h1 : _GEN_4610;
  assign _GEN_4612 = 9'h3a == _T_82861 ? 1'h1 : _GEN_4611;
  assign _GEN_4613 = 9'h3b == _T_82861 ? 1'h1 : _GEN_4612;
  assign _GEN_4614 = 9'h3c == _T_82861 ? 1'h1 : _GEN_4613;
  assign _GEN_4615 = 9'h3d == _T_82861 ? 1'h1 : _GEN_4614;
  assign _GEN_4616 = 9'h3e == _T_82861 ? 1'h1 : _GEN_4615;
  assign _GEN_4617 = 9'h3f == _T_82861 ? 1'h1 : _GEN_4616;
  assign _GEN_4618 = 9'h40 == _T_82861 ? _T_28219 : _GEN_4617;
  assign _GEN_4619 = 9'h41 == _T_82861 ? _T_27814 : _GEN_4618;
  assign _GEN_4620 = 9'h42 == _T_82861 ? _T_28597 : _GEN_4619;
  assign _GEN_4621 = 9'h43 == _T_82861 ? _T_28903 : _GEN_4620;
  assign _GEN_4622 = 9'h44 == _T_82861 ? 1'h1 : _GEN_4621;
  assign _GEN_4623 = 9'h45 == _T_82861 ? 1'h1 : _GEN_4622;
  assign _GEN_4624 = 9'h46 == _T_82861 ? 1'h1 : _GEN_4623;
  assign _GEN_4625 = 9'h47 == _T_82861 ? 1'h1 : _GEN_4624;
  assign _GEN_4626 = 9'h48 == _T_82861 ? 1'h1 : _GEN_4625;
  assign _GEN_4627 = 9'h49 == _T_82861 ? 1'h1 : _GEN_4626;
  assign _GEN_4628 = 9'h4a == _T_82861 ? 1'h1 : _GEN_4627;
  assign _GEN_4629 = 9'h4b == _T_82861 ? 1'h1 : _GEN_4628;
  assign _GEN_4630 = 9'h4c == _T_82861 ? 1'h1 : _GEN_4629;
  assign _GEN_4631 = 9'h4d == _T_82861 ? 1'h1 : _GEN_4630;
  assign _GEN_4632 = 9'h4e == _T_82861 ? 1'h1 : _GEN_4631;
  assign _GEN_4633 = 9'h4f == _T_82861 ? 1'h1 : _GEN_4632;
  assign _GEN_4634 = 9'h50 == _T_82861 ? 1'h1 : _GEN_4633;
  assign _GEN_4635 = 9'h51 == _T_82861 ? 1'h1 : _GEN_4634;
  assign _GEN_4636 = 9'h52 == _T_82861 ? 1'h1 : _GEN_4635;
  assign _GEN_4637 = 9'h53 == _T_82861 ? 1'h1 : _GEN_4636;
  assign _GEN_4638 = 9'h54 == _T_82861 ? 1'h1 : _GEN_4637;
  assign _GEN_4639 = 9'h55 == _T_82861 ? 1'h1 : _GEN_4638;
  assign _GEN_4640 = 9'h56 == _T_82861 ? 1'h1 : _GEN_4639;
  assign _GEN_4641 = 9'h57 == _T_82861 ? 1'h1 : _GEN_4640;
  assign _GEN_4642 = 9'h58 == _T_82861 ? 1'h1 : _GEN_4641;
  assign _GEN_4643 = 9'h59 == _T_82861 ? 1'h1 : _GEN_4642;
  assign _GEN_4644 = 9'h5a == _T_82861 ? 1'h1 : _GEN_4643;
  assign _GEN_4645 = 9'h5b == _T_82861 ? 1'h1 : _GEN_4644;
  assign _GEN_4646 = 9'h5c == _T_82861 ? 1'h1 : _GEN_4645;
  assign _GEN_4647 = 9'h5d == _T_82861 ? 1'h1 : _GEN_4646;
  assign _GEN_4648 = 9'h5e == _T_82861 ? 1'h1 : _GEN_4647;
  assign _GEN_4649 = 9'h5f == _T_82861 ? 1'h1 : _GEN_4648;
  assign _GEN_4650 = 9'h60 == _T_82861 ? 1'h1 : _GEN_4649;
  assign _GEN_4651 = 9'h61 == _T_82861 ? 1'h1 : _GEN_4650;
  assign _GEN_4652 = 9'h62 == _T_82861 ? 1'h1 : _GEN_4651;
  assign _GEN_4653 = 9'h63 == _T_82861 ? 1'h1 : _GEN_4652;
  assign _GEN_4654 = 9'h64 == _T_82861 ? 1'h1 : _GEN_4653;
  assign _GEN_4655 = 9'h65 == _T_82861 ? 1'h1 : _GEN_4654;
  assign _GEN_4656 = 9'h66 == _T_82861 ? 1'h1 : _GEN_4655;
  assign _GEN_4657 = 9'h67 == _T_82861 ? 1'h1 : _GEN_4656;
  assign _GEN_4658 = 9'h68 == _T_82861 ? 1'h1 : _GEN_4657;
  assign _GEN_4659 = 9'h69 == _T_82861 ? 1'h1 : _GEN_4658;
  assign _GEN_4660 = 9'h6a == _T_82861 ? 1'h1 : _GEN_4659;
  assign _GEN_4661 = 9'h6b == _T_82861 ? 1'h1 : _GEN_4660;
  assign _GEN_4662 = 9'h6c == _T_82861 ? 1'h1 : _GEN_4661;
  assign _GEN_4663 = 9'h6d == _T_82861 ? 1'h1 : _GEN_4662;
  assign _GEN_4664 = 9'h6e == _T_82861 ? 1'h1 : _GEN_4663;
  assign _GEN_4665 = 9'h6f == _T_82861 ? 1'h1 : _GEN_4664;
  assign _GEN_4666 = 9'h70 == _T_82861 ? 1'h1 : _GEN_4665;
  assign _GEN_4667 = 9'h71 == _T_82861 ? 1'h1 : _GEN_4666;
  assign _GEN_4668 = 9'h72 == _T_82861 ? 1'h1 : _GEN_4667;
  assign _GEN_4669 = 9'h73 == _T_82861 ? 1'h1 : _GEN_4668;
  assign _GEN_4670 = 9'h74 == _T_82861 ? 1'h1 : _GEN_4669;
  assign _GEN_4671 = 9'h75 == _T_82861 ? 1'h1 : _GEN_4670;
  assign _GEN_4672 = 9'h76 == _T_82861 ? 1'h1 : _GEN_4671;
  assign _GEN_4673 = 9'h77 == _T_82861 ? 1'h1 : _GEN_4672;
  assign _GEN_4674 = 9'h78 == _T_82861 ? 1'h1 : _GEN_4673;
  assign _GEN_4675 = 9'h79 == _T_82861 ? 1'h1 : _GEN_4674;
  assign _GEN_4676 = 9'h7a == _T_82861 ? 1'h1 : _GEN_4675;
  assign _GEN_4677 = 9'h7b == _T_82861 ? 1'h1 : _GEN_4676;
  assign _GEN_4678 = 9'h7c == _T_82861 ? 1'h1 : _GEN_4677;
  assign _GEN_4679 = 9'h7d == _T_82861 ? 1'h1 : _GEN_4678;
  assign _GEN_4680 = 9'h7e == _T_82861 ? 1'h1 : _GEN_4679;
  assign _GEN_4681 = 9'h7f == _T_82861 ? 1'h1 : _GEN_4680;
  assign _GEN_4682 = 9'h80 == _T_82861 ? 1'h1 : _GEN_4681;
  assign _GEN_4683 = 9'h81 == _T_82861 ? 1'h1 : _GEN_4682;
  assign _GEN_4684 = 9'h82 == _T_82861 ? 1'h1 : _GEN_4683;
  assign _GEN_4685 = 9'h83 == _T_82861 ? 1'h1 : _GEN_4684;
  assign _GEN_4686 = 9'h84 == _T_82861 ? 1'h1 : _GEN_4685;
  assign _GEN_4687 = 9'h85 == _T_82861 ? 1'h1 : _GEN_4686;
  assign _GEN_4688 = 9'h86 == _T_82861 ? 1'h1 : _GEN_4687;
  assign _GEN_4689 = 9'h87 == _T_82861 ? 1'h1 : _GEN_4688;
  assign _GEN_4690 = 9'h88 == _T_82861 ? 1'h1 : _GEN_4689;
  assign _GEN_4691 = 9'h89 == _T_82861 ? 1'h1 : _GEN_4690;
  assign _GEN_4692 = 9'h8a == _T_82861 ? 1'h1 : _GEN_4691;
  assign _GEN_4693 = 9'h8b == _T_82861 ? 1'h1 : _GEN_4692;
  assign _GEN_4694 = 9'h8c == _T_82861 ? 1'h1 : _GEN_4693;
  assign _GEN_4695 = 9'h8d == _T_82861 ? 1'h1 : _GEN_4694;
  assign _GEN_4696 = 9'h8e == _T_82861 ? 1'h1 : _GEN_4695;
  assign _GEN_4697 = 9'h8f == _T_82861 ? 1'h1 : _GEN_4696;
  assign _GEN_4698 = 9'h90 == _T_82861 ? 1'h1 : _GEN_4697;
  assign _GEN_4699 = 9'h91 == _T_82861 ? 1'h1 : _GEN_4698;
  assign _GEN_4700 = 9'h92 == _T_82861 ? 1'h1 : _GEN_4699;
  assign _GEN_4701 = 9'h93 == _T_82861 ? 1'h1 : _GEN_4700;
  assign _GEN_4702 = 9'h94 == _T_82861 ? 1'h1 : _GEN_4701;
  assign _GEN_4703 = 9'h95 == _T_82861 ? 1'h1 : _GEN_4702;
  assign _GEN_4704 = 9'h96 == _T_82861 ? 1'h1 : _GEN_4703;
  assign _GEN_4705 = 9'h97 == _T_82861 ? 1'h1 : _GEN_4704;
  assign _GEN_4706 = 9'h98 == _T_82861 ? 1'h1 : _GEN_4705;
  assign _GEN_4707 = 9'h99 == _T_82861 ? 1'h1 : _GEN_4706;
  assign _GEN_4708 = 9'h9a == _T_82861 ? 1'h1 : _GEN_4707;
  assign _GEN_4709 = 9'h9b == _T_82861 ? 1'h1 : _GEN_4708;
  assign _GEN_4710 = 9'h9c == _T_82861 ? 1'h1 : _GEN_4709;
  assign _GEN_4711 = 9'h9d == _T_82861 ? 1'h1 : _GEN_4710;
  assign _GEN_4712 = 9'h9e == _T_82861 ? 1'h1 : _GEN_4711;
  assign _GEN_4713 = 9'h9f == _T_82861 ? 1'h1 : _GEN_4712;
  assign _GEN_4714 = 9'ha0 == _T_82861 ? 1'h1 : _GEN_4713;
  assign _GEN_4715 = 9'ha1 == _T_82861 ? 1'h1 : _GEN_4714;
  assign _GEN_4716 = 9'ha2 == _T_82861 ? 1'h1 : _GEN_4715;
  assign _GEN_4717 = 9'ha3 == _T_82861 ? 1'h1 : _GEN_4716;
  assign _GEN_4718 = 9'ha4 == _T_82861 ? 1'h1 : _GEN_4717;
  assign _GEN_4719 = 9'ha5 == _T_82861 ? 1'h1 : _GEN_4718;
  assign _GEN_4720 = 9'ha6 == _T_82861 ? 1'h1 : _GEN_4719;
  assign _GEN_4721 = 9'ha7 == _T_82861 ? 1'h1 : _GEN_4720;
  assign _GEN_4722 = 9'ha8 == _T_82861 ? 1'h1 : _GEN_4721;
  assign _GEN_4723 = 9'ha9 == _T_82861 ? 1'h1 : _GEN_4722;
  assign _GEN_4724 = 9'haa == _T_82861 ? 1'h1 : _GEN_4723;
  assign _GEN_4725 = 9'hab == _T_82861 ? 1'h1 : _GEN_4724;
  assign _GEN_4726 = 9'hac == _T_82861 ? 1'h1 : _GEN_4725;
  assign _GEN_4727 = 9'had == _T_82861 ? 1'h1 : _GEN_4726;
  assign _GEN_4728 = 9'hae == _T_82861 ? 1'h1 : _GEN_4727;
  assign _GEN_4729 = 9'haf == _T_82861 ? 1'h1 : _GEN_4728;
  assign _GEN_4730 = 9'hb0 == _T_82861 ? 1'h1 : _GEN_4729;
  assign _GEN_4731 = 9'hb1 == _T_82861 ? 1'h1 : _GEN_4730;
  assign _GEN_4732 = 9'hb2 == _T_82861 ? 1'h1 : _GEN_4731;
  assign _GEN_4733 = 9'hb3 == _T_82861 ? 1'h1 : _GEN_4732;
  assign _GEN_4734 = 9'hb4 == _T_82861 ? 1'h1 : _GEN_4733;
  assign _GEN_4735 = 9'hb5 == _T_82861 ? 1'h1 : _GEN_4734;
  assign _GEN_4736 = 9'hb6 == _T_82861 ? 1'h1 : _GEN_4735;
  assign _GEN_4737 = 9'hb7 == _T_82861 ? 1'h1 : _GEN_4736;
  assign _GEN_4738 = 9'hb8 == _T_82861 ? 1'h1 : _GEN_4737;
  assign _GEN_4739 = 9'hb9 == _T_82861 ? 1'h1 : _GEN_4738;
  assign _GEN_4740 = 9'hba == _T_82861 ? 1'h1 : _GEN_4739;
  assign _GEN_4741 = 9'hbb == _T_82861 ? 1'h1 : _GEN_4740;
  assign _GEN_4742 = 9'hbc == _T_82861 ? 1'h1 : _GEN_4741;
  assign _GEN_4743 = 9'hbd == _T_82861 ? 1'h1 : _GEN_4742;
  assign _GEN_4744 = 9'hbe == _T_82861 ? 1'h1 : _GEN_4743;
  assign _GEN_4745 = 9'hbf == _T_82861 ? 1'h1 : _GEN_4744;
  assign _GEN_4746 = 9'hc0 == _T_82861 ? _T_27751 : _GEN_4745;
  assign _GEN_4747 = 9'hc1 == _T_82861 ? 1'h1 : _GEN_4746;
  assign _GEN_4748 = 9'hc2 == _T_82861 ? 1'h1 : _GEN_4747;
  assign _GEN_4749 = 9'hc3 == _T_82861 ? 1'h1 : _GEN_4748;
  assign _GEN_4750 = 9'hc4 == _T_82861 ? 1'h1 : _GEN_4749;
  assign _GEN_4751 = 9'hc5 == _T_82861 ? 1'h1 : _GEN_4750;
  assign _GEN_4752 = 9'hc6 == _T_82861 ? 1'h1 : _GEN_4751;
  assign _GEN_4753 = 9'hc7 == _T_82861 ? 1'h1 : _GEN_4752;
  assign _GEN_4754 = 9'hc8 == _T_82861 ? 1'h1 : _GEN_4753;
  assign _GEN_4755 = 9'hc9 == _T_82861 ? 1'h1 : _GEN_4754;
  assign _GEN_4756 = 9'hca == _T_82861 ? 1'h1 : _GEN_4755;
  assign _GEN_4757 = 9'hcb == _T_82861 ? 1'h1 : _GEN_4756;
  assign _GEN_4758 = 9'hcc == _T_82861 ? 1'h1 : _GEN_4757;
  assign _GEN_4759 = 9'hcd == _T_82861 ? 1'h1 : _GEN_4758;
  assign _GEN_4760 = 9'hce == _T_82861 ? _T_27571 : _GEN_4759;
  assign _GEN_4761 = 9'hcf == _T_82861 ? _T_29209 : _GEN_4760;
  assign _GEN_4762 = 9'hd0 == _T_82861 ? _T_28498 : _GEN_4761;
  assign _GEN_4763 = 9'hd1 == _T_82861 ? _T_28777 : _GEN_4762;
  assign _GEN_4764 = 9'hd2 == _T_82861 ? _T_29371 : _GEN_4763;
  assign _GEN_4765 = 9'hd3 == _T_82861 ? _T_27409 : _GEN_4764;
  assign _GEN_4766 = 9'hd4 == _T_82861 ? _T_28039 : _GEN_4765;
  assign _GEN_4767 = 9'hd5 == _T_82861 ? _T_28570 : _GEN_4766;
  assign _GEN_4768 = 9'hd6 == _T_82861 ? _T_29254 : _GEN_4767;
  assign _GEN_4769 = 9'hd7 == _T_82861 ? _T_29632 : _GEN_4768;
  assign _GEN_4770 = 9'hd8 == _T_82861 ? _T_27355 : _GEN_4769;
  assign _GEN_4771 = 9'hd9 == _T_82861 ? _T_27040 : _GEN_4770;
  assign _GEN_4772 = 9'hda == _T_82861 ? _T_29083 : _GEN_4771;
  assign _GEN_4773 = 9'hdb == _T_82861 ? _T_28399 : _GEN_4772;
  assign _GEN_4774 = 9'hdc == _T_82861 ? _T_27661 : _GEN_4773;
  assign _GEN_4775 = 9'hdd == _T_82861 ? _T_27481 : _GEN_4774;
  assign _GEN_4776 = 9'hde == _T_82861 ? _T_29650 : _GEN_4775;
  assign _GEN_4777 = 9'hdf == _T_82861 ? _T_28660 : _GEN_4776;
  assign _GEN_4778 = 9'he0 == _T_82861 ? _T_27895 : _GEN_4777;
  assign _GEN_4779 = 9'he1 == _T_82861 ? 1'h1 : _GEN_4778;
  assign _GEN_4780 = 9'he2 == _T_82861 ? 1'h1 : _GEN_4779;
  assign _GEN_4781 = 9'he3 == _T_82861 ? 1'h1 : _GEN_4780;
  assign _GEN_4782 = 9'he4 == _T_82861 ? 1'h1 : _GEN_4781;
  assign _GEN_4783 = 9'he5 == _T_82861 ? 1'h1 : _GEN_4782;
  assign _GEN_4784 = 9'he6 == _T_82861 ? 1'h1 : _GEN_4783;
  assign _GEN_4785 = 9'he7 == _T_82861 ? 1'h1 : _GEN_4784;
  assign _GEN_4786 = 9'he8 == _T_82861 ? 1'h1 : _GEN_4785;
  assign _GEN_4787 = 9'he9 == _T_82861 ? 1'h1 : _GEN_4786;
  assign _GEN_4788 = 9'hea == _T_82861 ? 1'h1 : _GEN_4787;
  assign _GEN_4789 = 9'heb == _T_82861 ? 1'h1 : _GEN_4788;
  assign _GEN_4790 = 9'hec == _T_82861 ? 1'h1 : _GEN_4789;
  assign _GEN_4791 = 9'hed == _T_82861 ? 1'h1 : _GEN_4790;
  assign _GEN_4792 = 9'hee == _T_82861 ? 1'h1 : _GEN_4791;
  assign _GEN_4793 = 9'hef == _T_82861 ? 1'h1 : _GEN_4792;
  assign _GEN_4794 = 9'hf0 == _T_82861 ? 1'h1 : _GEN_4793;
  assign _GEN_4795 = 9'hf1 == _T_82861 ? 1'h1 : _GEN_4794;
  assign _GEN_4796 = 9'hf2 == _T_82861 ? 1'h1 : _GEN_4795;
  assign _GEN_4797 = 9'hf3 == _T_82861 ? 1'h1 : _GEN_4796;
  assign _GEN_4798 = 9'hf4 == _T_82861 ? 1'h1 : _GEN_4797;
  assign _GEN_4799 = 9'hf5 == _T_82861 ? 1'h1 : _GEN_4798;
  assign _GEN_4800 = 9'hf6 == _T_82861 ? 1'h1 : _GEN_4799;
  assign _GEN_4801 = 9'hf7 == _T_82861 ? 1'h1 : _GEN_4800;
  assign _GEN_4802 = 9'hf8 == _T_82861 ? 1'h1 : _GEN_4801;
  assign _GEN_4803 = 9'hf9 == _T_82861 ? 1'h1 : _GEN_4802;
  assign _GEN_4804 = 9'hfa == _T_82861 ? 1'h1 : _GEN_4803;
  assign _GEN_4805 = 9'hfb == _T_82861 ? 1'h1 : _GEN_4804;
  assign _GEN_4806 = 9'hfc == _T_82861 ? 1'h1 : _GEN_4805;
  assign _GEN_4807 = 9'hfd == _T_82861 ? 1'h1 : _GEN_4806;
  assign _GEN_4808 = 9'hfe == _T_82861 ? 1'h1 : _GEN_4807;
  assign _GEN_4809 = 9'hff == _T_82861 ? 1'h1 : _GEN_4808;
  assign _GEN_4810 = 9'h100 == _T_82861 ? _T_27985 : _GEN_4809;
  assign _GEN_4811 = 9'h101 == _T_82861 ? _T_27220 : _GEN_4810;
  assign _GEN_4812 = 9'h102 == _T_82861 ? _T_29128 : _GEN_4811;
  assign _GEN_4813 = 9'h103 == _T_82861 ? _T_28300 : _GEN_4812;
  assign _GEN_4814 = 9'h104 == _T_82861 ? _T_27706 : _GEN_4813;
  assign _GEN_4815 = 9'h105 == _T_82861 ? _T_27346 : _GEN_4814;
  assign _GEN_4816 = 9'h106 == _T_82861 ? _T_29317 : _GEN_4815;
  assign _GEN_4817 = 9'h107 == _T_82861 ? _T_28885 : _GEN_4816;
  assign _GEN_4818 = 9'h108 == _T_82861 ? _T_28201 : _GEN_4817;
  assign _GEN_4819 = 9'h109 == _T_82861 ? _T_27535 : _GEN_4818;
  assign _GEN_4820 = 9'h10a == _T_82861 ? _T_28102 : _GEN_4819;
  assign _GEN_4821 = 9'h10b == _T_82861 ? _T_28696 : _GEN_4820;
  assign _GEN_4822 = 9'h10c == _T_82861 ? _T_29416 : _GEN_4821;
  assign _GEN_4823 = 9'h10d == _T_82861 ? _T_27103 : _GEN_4822;
  assign _GEN_4824 = 9'h10e == _T_82861 ? _T_27634 : _GEN_4823;
  assign _GEN_4825 = 9'h10f == _T_82861 ? _T_28489 : _GEN_4824;
  assign _GEN_4826 = 9'h110 == _T_82861 ? _T_29227 : _GEN_4825;
  assign _GEN_4827 = 9'h111 == _T_82861 ? _T_29344 : _GEN_4826;
  assign _GEN_4828 = 9'h112 == _T_82861 ? _T_28408 : _GEN_4827;
  assign _GEN_4829 = 9'h113 == _T_82861 ? _T_27778 : _GEN_4828;
  assign _GEN_4830 = 9'h114 == _T_82861 ? _T_27049 : _GEN_4829;
  assign _GEN_4831 = 9'h115 == _T_82861 ? _T_29542 : _GEN_4830;
  assign _GEN_4832 = 9'h116 == _T_82861 ? _T_28642 : _GEN_4831;
  assign _GEN_4833 = 9'h117 == _T_82861 ? _T_28210 : _GEN_4832;
  assign _GEN_4834 = 9'h118 == _T_82861 ? _T_27472 : _GEN_4833;
  assign _GEN_4835 = 9'h119 == _T_82861 ? _T_28291 : _GEN_4834;
  assign _GEN_4836 = 9'h11a == _T_82861 ? _T_28849 : _GEN_4835;
  assign _GEN_4837 = 9'h11b == _T_82861 ? _T_29470 : _GEN_4836;
  assign _GEN_4838 = 9'h11c == _T_82861 ? _T_27292 : _GEN_4837;
  assign _GEN_4839 = 9'h11d == _T_82861 ? _T_27886 : _GEN_4838;
  assign _GEN_4840 = 9'h11e == _T_82861 ? _T_28273 : _GEN_4839;
  assign _GEN_4841 = 9'h11f == _T_82861 ? _T_29263 : _GEN_4840;
  assign _GEN_4842 = 9'h120 == _T_82861 ? _T_27184 : _GEN_4841;
  assign _GEN_4843 = 9'h121 == _T_82861 ? _T_27319 : _GEN_4842;
  assign _GEN_4844 = 9'h122 == _T_82861 ? _T_29173 : _GEN_4843;
  assign _GEN_4845 = 9'h123 == _T_82861 ? _T_28282 : _GEN_4844;
  assign _GEN_4846 = 9'h124 == _T_82861 ? _T_27589 : _GEN_4845;
  assign _GEN_4847 = 9'h125 == _T_82861 ? _T_27490 : _GEN_4846;
  assign _GEN_4848 = 9'h126 == _T_82861 ? _T_29389 : _GEN_4847;
  assign _GEN_4849 = 9'h127 == _T_82861 ? _T_28840 : _GEN_4848;
  assign _GEN_4850 = 9'h128 == _T_82861 ? _T_28228 : _GEN_4849;
  assign _GEN_4851 = 9'h129 == _T_82861 ? _T_27733 : _GEN_4850;
  assign _GEN_4852 = 9'h12a == _T_82861 ? _T_28156 : _GEN_4851;
  assign _GEN_4853 = 9'h12b == _T_82861 ? _T_28687 : _GEN_4852;
  assign _GEN_4854 = 9'h12c == _T_82861 ? _T_29272 : _GEN_4853;
  assign _GEN_4855 = 9'h12d == _T_82861 ? _T_27193 : _GEN_4854;
  assign _GEN_4856 = 9'h12e == _T_82861 ? _T_27697 : _GEN_4855;
  assign _GEN_4857 = 9'h12f == _T_82861 ? _T_28480 : _GEN_4856;
  assign _GEN_4858 = 9'h130 == _T_82861 ? _T_29119 : _GEN_4857;
  assign _GEN_4859 = 9'h131 == _T_82861 ? _T_29362 : _GEN_4858;
  assign _GEN_4860 = 9'h132 == _T_82861 ? _T_28678 : _GEN_4859;
  assign _GEN_4861 = 9'h133 == _T_82861 ? _T_27580 : _GEN_4860;
  assign _GEN_4862 = 9'h134 == _T_82861 ? _T_27058 : _GEN_4861;
  assign _GEN_4863 = 9'h135 == _T_82861 ? _T_29623 : _GEN_4862;
  assign _GEN_4864 = 9'h136 == _T_82861 ? _T_28894 : _GEN_4863;
  assign _GEN_4865 = 9'h137 == _T_82861 ? _T_28129 : _GEN_4864;
  assign _GEN_4866 = 9'h138 == _T_82861 ? _T_27562 : _GEN_4865;
  assign _GEN_4867 = 9'h139 == _T_82861 ? _T_28345 : _GEN_4866;
  assign _GEN_4868 = 9'h13a == _T_82861 ? _T_29002 : _GEN_4867;
  assign _GEN_4869 = 9'h13b == _T_82861 ? _T_29290 : _GEN_4868;
  assign _GEN_4870 = 9'h13c == _T_82861 ? _T_27337 : _GEN_4869;
  assign _GEN_4871 = 9'h13d == _T_82861 ? _T_27913 : _GEN_4870;
  assign _GEN_4872 = 9'h13e == _T_82861 ? _T_28453 : _GEN_4871;
  assign _GEN_4873 = 9'h13f == _T_82861 ? _T_29110 : _GEN_4872;
  assign _GEN_4874 = 9'h140 == _T_82861 ? _T_27202 : _GEN_4873;
  assign _GEN_4875 = 9'h141 == _T_82861 ? _T_27391 : _GEN_4874;
  assign _GEN_4876 = 9'h142 == _T_82861 ? _T_29578 : _GEN_4875;
  assign _GEN_4877 = 9'h143 == _T_82861 ? _T_28561 : _GEN_4876;
  assign _GEN_4878 = 9'h144 == _T_82861 ? _T_27877 : _GEN_4877;
  assign _GEN_4879 = 9'h145 == _T_82861 ? _T_27310 : _GEN_4878;
  assign _GEN_4880 = 9'h146 == _T_82861 ? _T_29380 : _GEN_4879;
  assign _GEN_4881 = 9'h147 == _T_82861 ? _T_28867 : _GEN_4880;
  assign _GEN_4882 = 9'h148 == _T_82861 ? _T_27967 : _GEN_4881;
  assign _GEN_4883 = 9'h149 == _T_82861 ? _T_27832 : _GEN_4882;
  assign _GEN_4884 = 9'h14a == _T_82861 ? _T_28606 : _GEN_4883;
  assign _GEN_4885 = 9'h14b == _T_82861 ? _T_28912 : _GEN_4884;
  assign _GEN_4886 = 9'h14c == _T_82861 ? _T_29506 : _GEN_4885;
  assign _GEN_4887 = 9'h14d == _T_82861 ? _T_26977 : _GEN_4886;
  assign _GEN_4888 = 9'h14e == _T_82861 ? _T_27688 : _GEN_4887;
  assign _GEN_4889 = 9'h14f == _T_82861 ? _T_28372 : _GEN_4888;
  assign _GEN_4890 = 9'h150 == _T_82861 ? _T_28984 : _GEN_4889;
  assign _GEN_4891 = 9'h151 == _T_82861 ? _T_29596 : _GEN_4890;
  assign _GEN_4892 = 9'h152 == _T_82861 ? _T_28957 : _GEN_4891;
  assign _GEN_4893 = 9'h153 == _T_82861 ? _T_28003 : _GEN_4892;
  assign _GEN_4894 = 9'h154 == _T_82861 ? _T_27157 : _GEN_4893;
  assign _GEN_4895 = 9'h155 == _T_82861 ? _T_29398 : _GEN_4894;
  assign _GEN_4896 = 9'h156 == _T_82861 ? _T_28804 : _GEN_4895;
  assign _GEN_4897 = 9'h157 == _T_82861 ? _T_28093 : _GEN_4896;
  assign _GEN_4898 = 9'h158 == _T_82861 ? _T_27256 : _GEN_4897;
  assign _GEN_4899 = 9'h159 == _T_82861 ? _T_28534 : _GEN_4898;
  assign _GEN_4900 = 9'h15a == _T_82861 ? _T_29245 : _GEN_4899;
  assign _GEN_4901 = 9'h15b == _T_82861 ? _T_26968 : _GEN_4900;
  assign _GEN_4902 = 9'h15c == _T_82861 ? _T_27436 : _GEN_4901;
  assign _GEN_4903 = 9'h15d == _T_82861 ? _T_27715 : _GEN_4902;
  assign _GEN_4904 = 9'h15e == _T_82861 ? _T_28381 : _GEN_4903;
  assign _GEN_4905 = 9'h15f == _T_82861 ? _T_29137 : _GEN_4904;
  assign _GEN_4906 = 9'h160 == _T_82861 ? _T_27013 : _GEN_4905;
  assign _GEN_4907 = 9'h161 == _T_82861 ? _T_27445 : _GEN_4906;
  assign _GEN_4908 = 9'h162 == _T_82861 ? _T_29614 : _GEN_4907;
  assign _GEN_4909 = 9'h163 == _T_82861 ? _T_28813 : _GEN_4908;
  assign _GEN_4910 = 9'h164 == _T_82861 ? _T_27940 : _GEN_4909;
  assign _GEN_4911 = 9'h165 == _T_82861 ? _T_27265 : _GEN_4910;
  assign _GEN_4912 = 9'h166 == _T_82861 ? _T_29425 : _GEN_4911;
  assign _GEN_4913 = 9'h167 == _T_82861 ? _T_28975 : _GEN_4912;
  assign _GEN_4914 = 9'h168 == _T_82861 ? _T_28111 : _GEN_4913;
  assign _GEN_4915 = 9'h169 == _T_82861 ? _T_27805 : _GEN_4914;
  assign _GEN_4916 = 9'h16a == _T_82861 ? _T_28435 : _GEN_4915;
  assign _GEN_4917 = 9'h16b == _T_82861 ? _T_29047 : _GEN_4916;
  assign _GEN_4918 = 9'h16c == _T_82861 ? _T_29677 : _GEN_4917;
  assign _GEN_4919 = 9'h16d == _T_82861 ? _T_26950 : _GEN_4918;
  assign _GEN_4920 = 9'h16e == _T_82861 ? _T_27670 : _GEN_4919;
  assign _GEN_4921 = 9'h16f == _T_82861 ? _T_28543 : _GEN_4920;
  assign _GEN_4922 = 9'h170 == _T_82861 ? _T_29092 : _GEN_4921;
  assign _GEN_4923 = 9'h171 == _T_82861 ? _T_29569 : _GEN_4922;
  assign _GEN_4924 = 9'h172 == _T_82861 ? _T_28930 : _GEN_4923;
  assign _GEN_4925 = 9'h173 == _T_82861 ? _T_28075 : _GEN_4924;
  assign _GEN_4926 = 9'h174 == _T_82861 ? _T_27238 : _GEN_4925;
  assign _GEN_4927 = 9'h175 == _T_82861 ? _T_29353 : _GEN_4926;
  assign _GEN_4928 = 9'h176 == _T_82861 ? _T_28768 : _GEN_4927;
  assign _GEN_4929 = 9'h177 == _T_82861 ? _T_28246 : _GEN_4928;
  assign _GEN_4930 = 9'h178 == _T_82861 ? _T_27400 : _GEN_4929;
  assign _GEN_4931 = 9'h179 == _T_82861 ? _T_28426 : _GEN_4930;
  assign _GEN_4932 = 9'h17a == _T_82861 ? _T_29182 : _GEN_4931;
  assign _GEN_4933 = 9'h17b == _T_82861 ? _T_27076 : _GEN_4932;
  assign _GEN_4934 = 9'h17c == _T_82861 ? _T_27607 : _GEN_4933;
  assign _GEN_4935 = 9'h17d == _T_82861 ? _T_27652 : _GEN_4934;
  assign _GEN_4936 = 9'h17e == _T_82861 ? _T_28336 : _GEN_4935;
  assign _GEN_4937 = 9'h17f == _T_82861 ? _T_29236 : _GEN_4936;
  assign _GEN_4938 = 9'h180 == _T_82861 ? _T_27121 : _GEN_4937;
  assign _GEN_4939 = 9'h181 == _T_82861 ? _T_27112 : _GEN_4938;
  assign _GEN_4940 = 9'h182 == _T_82861 ? _T_28993 : _GEN_4939;
  assign _GEN_4941 = 9'h183 == _T_82861 ? _T_28516 : _GEN_4940;
  assign _GEN_4942 = 9'h184 == _T_82861 ? _T_27931 : _GEN_4941;
  assign _GEN_4943 = 9'h185 == _T_82861 ? _T_27229 : _GEN_4942;
  assign _GEN_4944 = 9'h186 == _T_82861 ? _T_29146 : _GEN_4943;
  assign _GEN_4945 = 9'h187 == _T_82861 ? _T_28318 : _GEN_4944;
  assign _GEN_4946 = 9'h188 == _T_82861 ? _T_27724 : _GEN_4945;
  assign _GEN_4947 = 9'h189 == _T_82861 ? _T_28048 : _GEN_4946;
  assign _GEN_4948 = 9'h18a == _T_82861 ? _T_28669 : _GEN_4947;
  assign _GEN_4949 = 9'h18b == _T_82861 ? _T_29488 : _GEN_4948;
  assign _GEN_4950 = 9'h18c == _T_82861 ? _T_27508 : _GEN_4949;
  assign _GEN_4951 = 9'h18d == _T_82861 ? _T_27463 : _GEN_4950;
  assign _GEN_4952 = 9'h18e == _T_82861 ? _T_28138 : _GEN_4951;
  assign _GEN_4953 = 9'h18f == _T_82861 ? _T_28633 : _GEN_4952;
  assign _GEN_4954 = 9'h190 == _T_82861 ? _T_29452 : _GEN_4953;
  assign _GEN_4955 = 9'h191 == _T_82861 ? _T_29155 : _GEN_4954;
  assign _GEN_4956 = 9'h192 == _T_82861 ? _T_28264 : _GEN_4955;
  assign _GEN_4957 = 9'h193 == _T_82861 ? _T_27922 : _GEN_4956;
  assign _GEN_4958 = 9'h194 == _T_82861 ? _T_27166 : _GEN_4957;
  assign _GEN_4959 = 9'h195 == _T_82861 ? _T_29326 : _GEN_4958;
  assign _GEN_4960 = 9'h196 == _T_82861 ? _T_28390 : _GEN_4959;
  assign _GEN_4961 = 9'h197 == _T_82861 ? _T_27760 : _GEN_4960;
  assign _GEN_4962 = 9'h198 == _T_82861 ? _T_27022 : _GEN_4961;
  assign _GEN_4963 = 9'h199 == _T_82861 ? _T_28876 : _GEN_4962;
  assign _GEN_4964 = 9'h19a == _T_82861 ? _T_29308 : _GEN_4963;
  assign _GEN_4965 = 9'h19b == _T_82861 ? _T_27517 : _GEN_4964;
  assign _GEN_4966 = 9'h19c == _T_82861 ? _T_28165 : _GEN_4965;
  assign _GEN_4967 = 9'h19d == _T_82861 ? _T_28309 : _GEN_4966;
  assign _GEN_4968 = 9'h19e == _T_82861 ? _T_28858 : _GEN_4967;
  assign _GEN_4969 = 9'h19f == _T_82861 ? _T_29479 : _GEN_4968;
  assign _GEN_4970 = 9'h1a0 == _T_82861 ? _T_27301 : _GEN_4969;
  assign _GEN_4971 = 9'h1a1 == _T_82861 ? _T_27175 : _GEN_4970;
  assign _GEN_4972 = 9'h1a2 == _T_82861 ? _T_29164 : _GEN_4971;
  assign _GEN_4973 = 9'h1a3 == _T_82861 ? _T_28417 : _GEN_4972;
  assign _GEN_4974 = 9'h1a4 == _T_82861 ? _T_27949 : _GEN_4973;
  assign _GEN_4975 = 9'h1a5 == _T_82861 ? _T_27283 : _GEN_4974;
  assign _GEN_4976 = 9'h1a6 == _T_82861 ? _T_29335 : _GEN_4975;
  assign _GEN_4977 = 9'h1a7 == _T_82861 ? _T_28255 : _GEN_4976;
  assign _GEN_4978 = 9'h1a8 == _T_82861 ? _T_27742 : _GEN_4977;
  assign _GEN_4979 = 9'h1a9 == _T_82861 ? _T_28174 : _GEN_4978;
  assign _GEN_4980 = 9'h1aa == _T_82861 ? _T_28750 : _GEN_4979;
  assign _GEN_4981 = 9'h1ab == _T_82861 ? _T_29515 : _GEN_4980;
  assign _GEN_4982 = 9'h1ac == _T_82861 ? _T_27526 : _GEN_4981;
  assign _GEN_4983 = 9'h1ad == _T_82861 ? _T_27769 : _GEN_4982;
  assign _GEN_4984 = 9'h1ae == _T_82861 ? _T_28192 : _GEN_4983;
  assign _GEN_4985 = 9'h1af == _T_82861 ? _T_28723 : _GEN_4984;
  assign _GEN_4986 = 9'h1b0 == _T_82861 ? _T_29299 : _GEN_4985;
  assign _GEN_4987 = 9'h1b1 == _T_82861 ? _T_29191 : _GEN_4986;
  assign _GEN_4988 = 9'h1b2 == _T_82861 ? _T_28471 : _GEN_4987;
  assign _GEN_4989 = 9'h1b3 == _T_82861 ? _T_27823 : _GEN_4988;
  assign _GEN_4990 = 9'h1b4 == _T_82861 ? _T_27211 : _GEN_4989;
  assign _GEN_4991 = 9'h1b5 == _T_82861 ? _T_29434 : _GEN_4990;
  assign _GEN_4992 = 9'h1b6 == _T_82861 ? _T_28714 : _GEN_4991;
  assign _GEN_4993 = 9'h1b7 == _T_82861 ? _T_27625 : _GEN_4992;
  assign _GEN_4994 = 9'h1b8 == _T_82861 ? _T_27085 : _GEN_4993;
  assign _GEN_4995 = 9'h1b9 == _T_82861 ? _T_28921 : _GEN_4994;
  assign _GEN_4996 = 9'h1ba == _T_82861 ? _T_29551 : _GEN_4995;
  assign _GEN_4997 = 9'h1bb == _T_82861 ? _T_27382 : _GEN_4996;
  assign _GEN_4998 = 9'h1bc == _T_82861 ? _T_28237 : _GEN_4997;
  assign _GEN_4999 = 9'h1bd == _T_82861 ? _T_28327 : _GEN_4998;
  assign _GEN_5000 = 9'h1be == _T_82861 ? _T_29011 : _GEN_4999;
  assign _GEN_5001 = 9'h1bf == _T_82861 ? _T_29281 : _GEN_5000;
  assign _GEN_5002 = 9'h1c0 == _T_82861 ? _T_27328 : _GEN_5001;
  assign _GEN_5003 = 9'h1c1 == _T_82861 ? _T_27067 : _GEN_5002;
  assign _GEN_5004 = 9'h1c2 == _T_82861 ? _T_29038 : _GEN_5003;
  assign _GEN_5005 = 9'h1c3 == _T_82861 ? _T_28444 : _GEN_5004;
  assign _GEN_5006 = 9'h1c4 == _T_82861 ? _T_27598 : _GEN_5005;
  assign _GEN_5007 = 9'h1c5 == _T_82861 ? _T_27499 : _GEN_5006;
  assign _GEN_5008 = 9'h1c6 == _T_82861 ? _T_29668 : _GEN_5007;
  assign _GEN_5009 = 9'h1c7 == _T_82861 ? _T_28651 : _GEN_5008;
  assign _GEN_5010 = 9'h1c8 == _T_82861 ? _T_27868 : _GEN_5009;
  assign _GEN_5011 = 9'h1c9 == _T_82861 ? _T_28066 : _GEN_5010;
  assign _GEN_5012 = 9'h1ca == _T_82861 ? _T_28822 : _GEN_5011;
  assign _GEN_5013 = 9'h1cb == _T_82861 ? _T_29533 : _GEN_5012;
  assign _GEN_5014 = 9'h1cc == _T_82861 ? _T_27274 : _GEN_5013;
  assign _GEN_5015 = 9'h1cd == _T_82861 ? _T_27850 : _GEN_5014;
  assign _GEN_5016 = 9'h1ce == _T_82861 ? _T_28615 : _GEN_5015;
  assign _GEN_5017 = 9'h1cf == _T_82861 ? _T_28948 : _GEN_5016;
  assign _GEN_5018 = 9'h1d0 == _T_82861 ? _T_29497 : _GEN_5017;
  assign _GEN_5019 = 9'h1d1 == _T_82861 ? _T_29029 : _GEN_5018;
  assign _GEN_5020 = 9'h1d2 == _T_82861 ? _T_28363 : _GEN_5019;
  assign _GEN_5021 = 9'h1d3 == _T_82861 ? _T_27787 : _GEN_5020;
  assign _GEN_5022 = 9'h1d4 == _T_82861 ? _T_26995 : _GEN_5021;
  assign _GEN_5023 = 9'h1d5 == _T_82861 ? _T_29605 : _GEN_5022;
  assign _GEN_5024 = 9'h1d6 == _T_82861 ? _T_28966 : _GEN_5023;
  assign _GEN_5025 = 9'h1d7 == _T_82861 ? _T_27976 : _GEN_5024;
  assign _GEN_5026 = 9'h1d8 == _T_82861 ? _T_27148 : _GEN_5025;
  assign _GEN_5027 = 9'h1d9 == _T_82861 ? _T_28732 : _GEN_5026;
  assign _GEN_5028 = 9'h1da == _T_82861 ? _T_29443 : _GEN_5027;
  assign _GEN_5029 = 9'h1db == _T_82861 ? _T_27364 : _GEN_5028;
  assign _GEN_5030 = 9'h1dc == _T_82861 ? _T_28012 : _GEN_5029;
  assign _GEN_5031 = 9'h1dd == _T_82861 ? _T_28507 : _GEN_5030;
  assign _GEN_5032 = 9'h1de == _T_82861 ? _T_29218 : _GEN_5031;
  assign _GEN_5033 = 9'h1df == _T_82861 ? _T_26959 : _GEN_5032;
  assign _GEN_5034 = 9'h1e0 == _T_82861 ? _T_27454 : _GEN_5033;
  assign _GEN_5035 = 9'h1e1 == _T_82861 ? _T_27004 : _GEN_5034;
  assign _GEN_5036 = 9'h1e2 == _T_82861 ? _T_29056 : _GEN_5035;
  assign _GEN_5037 = 9'h1e3 == _T_82861 ? _T_28579 : _GEN_5036;
  assign _GEN_5038 = 9'h1e4 == _T_82861 ? _T_27796 : _GEN_5037;
  assign _GEN_5039 = 9'h1e5 == _T_82861 ? _T_27418 : _GEN_5038;
  assign _GEN_5040 = 9'h1e6 == _T_82861 ? _T_29587 : _GEN_5039;
  assign _GEN_5041 = 9'h1e7 == _T_82861 ? _T_28786 : _GEN_5040;
  assign _GEN_5042 = 9'h1e8 == _T_82861 ? _T_27994 : _GEN_5041;
  assign _GEN_5043 = 9'h1e9 == _T_82861 ? _T_28030 : _GEN_5042;
  assign _GEN_5044 = 9'h1ea == _T_82861 ? _T_28741 : _GEN_5043;
  assign _GEN_5045 = 9'h1eb == _T_82861 ? _T_29641 : _GEN_5044;
  assign _GEN_5046 = 9'h1ec == _T_82861 ? _T_27373 : _GEN_5045;
  assign _GEN_5047 = 9'h1ed == _T_82861 ? _T_27859 : _GEN_5046;
  assign _GEN_5048 = 9'h1ee == _T_82861 ? _T_28525 : _GEN_5047;
  assign _GEN_5049 = 9'h1ef == _T_82861 ? _T_29074 : _GEN_5048;
  assign _GEN_5050 = 9'h1f0 == _T_82861 ? _T_29659 : _GEN_5049;
  assign _GEN_5051 = 9'h1f1 == _T_82861 ? _T_29020 : _GEN_5050;
  assign _GEN_5052 = 9'h1f2 == _T_82861 ? _T_28354 : _GEN_5051;
  assign _GEN_5053 = 9'h1f3 == _T_82861 ? _T_27958 : _GEN_5052;
  assign _GEN_5054 = 9'h1f4 == _T_82861 ? _T_27139 : _GEN_5053;
  assign _GEN_5055 = 9'h1f5 == _T_82861 ? _T_29560 : _GEN_5054;
  assign _GEN_5056 = 9'h1f6 == _T_82861 ? _T_28939 : _GEN_5055;
  assign _GEN_5057 = 9'h1f7 == _T_82861 ? _T_28084 : _GEN_5056;
  assign _GEN_5058 = 9'h1f8 == _T_82861 ? _T_27247 : _GEN_5057;
  assign _GEN_5059 = 9'h1f9 == _T_82861 ? _T_28705 : _GEN_5058;
  assign _GEN_5060 = 9'h1fa == _T_82861 ? _T_29407 : _GEN_5059;
  assign _GEN_5061 = 9'h1fb == _T_82861 ? _T_27544 : _GEN_5060;
  assign _GEN_5062 = 9'h1fc == _T_82861 ? _T_28120 : _GEN_5061;
  assign _GEN_5063 = 9'h1fd == _T_82861 ? _T_28462 : _GEN_5062;
  assign _GEN_5064 = 9'h1fe == _T_82861 ? _T_29200 : _GEN_5063;
  assign _GEN_5065 = 9'h1ff == _T_82861 ? _T_27094 : _GEN_5064;
  assign _GEN_5066 = 9'h1 == _T_82861 ? 32'h4c0006f : 32'hc0006f;
  assign _GEN_5067 = 9'h2 == _T_82861 ? 32'h340006f : _GEN_5066;
  assign _GEN_5068 = 9'h3 == _T_82861 ? 32'hff0000f : _GEN_5067;
  assign _GEN_5069 = 9'h4 == _T_82861 ? 32'h7b241073 : _GEN_5068;
  assign _GEN_5070 = 9'h5 == _T_82861 ? 32'hf1402473 : _GEN_5069;
  assign _GEN_5071 = 9'h6 == _T_82861 ? 32'h10802023 : _GEN_5070;
  assign _GEN_5072 = 9'h7 == _T_82861 ? 32'h40044403 : _GEN_5071;
  assign _GEN_5073 = 9'h8 == _T_82861 ? 32'h147413 : _GEN_5072;
  assign _GEN_5074 = 9'h9 == _T_82861 ? 32'h2041063 : _GEN_5073;
  assign _GEN_5075 = 9'ha == _T_82861 ? 32'hf1402473 : _GEN_5074;
  assign _GEN_5076 = 9'hb == _T_82861 ? 32'h40044403 : _GEN_5075;
  assign _GEN_5077 = 9'hc == _T_82861 ? 32'h247413 : _GEN_5076;
  assign _GEN_5078 = 9'hd == _T_82861 ? 32'hfc0418e3 : _GEN_5077;
  assign _GEN_5079 = 9'he == _T_82861 ? 32'hfddff06f : _GEN_5078;
  assign _GEN_5080 = 9'hf == _T_82861 ? 32'h10002623 : _GEN_5079;
  assign _GEN_5081 = 9'h10 == _T_82861 ? 32'h100073 : _GEN_5080;
  assign _GEN_5082 = 9'h11 == _T_82861 ? 32'h7b202473 : _GEN_5081;
  assign _GEN_5083 = 9'h12 == _T_82861 ? 32'h10002223 : _GEN_5082;
  assign _GEN_5084 = 9'h13 == _T_82861 ? 32'h30000067 : _GEN_5083;
  assign _GEN_5085 = 9'h14 == _T_82861 ? 32'hf1402473 : _GEN_5084;
  assign _GEN_5086 = 9'h15 == _T_82861 ? 32'h10802423 : _GEN_5085;
  assign _GEN_5087 = 9'h16 == _T_82861 ? 32'h7b202473 : _GEN_5086;
  assign _GEN_5088 = 9'h17 == _T_82861 ? 32'h7b200073 : _GEN_5087;
  assign _GEN_5089 = 9'h18 == _T_82861 ? 32'h0 : _GEN_5088;
  assign _GEN_5090 = 9'h19 == _T_82861 ? 32'h0 : _GEN_5089;
  assign _GEN_5091 = 9'h1a == _T_82861 ? 32'h0 : _GEN_5090;
  assign _GEN_5092 = 9'h1b == _T_82861 ? 32'h0 : _GEN_5091;
  assign _GEN_5093 = 9'h1c == _T_82861 ? 32'h0 : _GEN_5092;
  assign _GEN_5094 = 9'h1d == _T_82861 ? 32'h0 : _GEN_5093;
  assign _GEN_5095 = 9'h1e == _T_82861 ? 32'h0 : _GEN_5094;
  assign _GEN_5096 = 9'h1f == _T_82861 ? 32'h0 : _GEN_5095;
  assign _GEN_5097 = 9'h20 == _T_82861 ? 32'h0 : _GEN_5096;
  assign _GEN_5098 = 9'h21 == _T_82861 ? 32'h0 : _GEN_5097;
  assign _GEN_5099 = 9'h22 == _T_82861 ? 32'h0 : _GEN_5098;
  assign _GEN_5100 = 9'h23 == _T_82861 ? 32'h0 : _GEN_5099;
  assign _GEN_5101 = 9'h24 == _T_82861 ? 32'h0 : _GEN_5100;
  assign _GEN_5102 = 9'h25 == _T_82861 ? 32'h0 : _GEN_5101;
  assign _GEN_5103 = 9'h26 == _T_82861 ? 32'h0 : _GEN_5102;
  assign _GEN_5104 = 9'h27 == _T_82861 ? 32'h0 : _GEN_5103;
  assign _GEN_5105 = 9'h28 == _T_82861 ? 32'h0 : _GEN_5104;
  assign _GEN_5106 = 9'h29 == _T_82861 ? 32'h0 : _GEN_5105;
  assign _GEN_5107 = 9'h2a == _T_82861 ? 32'h0 : _GEN_5106;
  assign _GEN_5108 = 9'h2b == _T_82861 ? 32'h0 : _GEN_5107;
  assign _GEN_5109 = 9'h2c == _T_82861 ? 32'h0 : _GEN_5108;
  assign _GEN_5110 = 9'h2d == _T_82861 ? 32'h0 : _GEN_5109;
  assign _GEN_5111 = 9'h2e == _T_82861 ? 32'h0 : _GEN_5110;
  assign _GEN_5112 = 9'h2f == _T_82861 ? 32'h0 : _GEN_5111;
  assign _GEN_5113 = 9'h30 == _T_82861 ? 32'h0 : _GEN_5112;
  assign _GEN_5114 = 9'h31 == _T_82861 ? 32'h0 : _GEN_5113;
  assign _GEN_5115 = 9'h32 == _T_82861 ? 32'h0 : _GEN_5114;
  assign _GEN_5116 = 9'h33 == _T_82861 ? 32'h0 : _GEN_5115;
  assign _GEN_5117 = 9'h34 == _T_82861 ? 32'h0 : _GEN_5116;
  assign _GEN_5118 = 9'h35 == _T_82861 ? 32'h0 : _GEN_5117;
  assign _GEN_5119 = 9'h36 == _T_82861 ? 32'h0 : _GEN_5118;
  assign _GEN_5120 = 9'h37 == _T_82861 ? 32'h0 : _GEN_5119;
  assign _GEN_5121 = 9'h38 == _T_82861 ? 32'h0 : _GEN_5120;
  assign _GEN_5122 = 9'h39 == _T_82861 ? 32'h0 : _GEN_5121;
  assign _GEN_5123 = 9'h3a == _T_82861 ? 32'h0 : _GEN_5122;
  assign _GEN_5124 = 9'h3b == _T_82861 ? 32'h0 : _GEN_5123;
  assign _GEN_5125 = 9'h3c == _T_82861 ? 32'h0 : _GEN_5124;
  assign _GEN_5126 = 9'h3d == _T_82861 ? 32'h0 : _GEN_5125;
  assign _GEN_5127 = 9'h3e == _T_82861 ? 32'h0 : _GEN_5126;
  assign _GEN_5128 = 9'h3f == _T_82861 ? 32'h0 : _GEN_5127;
  assign _GEN_5129 = 9'h40 == _T_82861 ? _T_102902_64 : _GEN_5128;
  assign _GEN_5130 = 9'h41 == _T_82861 ? _T_102902_65 : _GEN_5129;
  assign _GEN_5131 = 9'h42 == _T_82861 ? _T_102902_66 : _GEN_5130;
  assign _GEN_5132 = 9'h43 == _T_82861 ? _T_102902_67 : _GEN_5131;
  assign _GEN_5133 = 9'h44 == _T_82861 ? 32'h0 : _GEN_5132;
  assign _GEN_5134 = 9'h45 == _T_82861 ? 32'h0 : _GEN_5133;
  assign _GEN_5135 = 9'h46 == _T_82861 ? 32'h0 : _GEN_5134;
  assign _GEN_5136 = 9'h47 == _T_82861 ? 32'h0 : _GEN_5135;
  assign _GEN_5137 = 9'h48 == _T_82861 ? 32'h0 : _GEN_5136;
  assign _GEN_5138 = 9'h49 == _T_82861 ? 32'h0 : _GEN_5137;
  assign _GEN_5139 = 9'h4a == _T_82861 ? 32'h0 : _GEN_5138;
  assign _GEN_5140 = 9'h4b == _T_82861 ? 32'h0 : _GEN_5139;
  assign _GEN_5141 = 9'h4c == _T_82861 ? 32'h0 : _GEN_5140;
  assign _GEN_5142 = 9'h4d == _T_82861 ? 32'h0 : _GEN_5141;
  assign _GEN_5143 = 9'h4e == _T_82861 ? 32'h0 : _GEN_5142;
  assign _GEN_5144 = 9'h4f == _T_82861 ? 32'h0 : _GEN_5143;
  assign _GEN_5145 = 9'h50 == _T_82861 ? 32'h0 : _GEN_5144;
  assign _GEN_5146 = 9'h51 == _T_82861 ? 32'h0 : _GEN_5145;
  assign _GEN_5147 = 9'h52 == _T_82861 ? 32'h0 : _GEN_5146;
  assign _GEN_5148 = 9'h53 == _T_82861 ? 32'h0 : _GEN_5147;
  assign _GEN_5149 = 9'h54 == _T_82861 ? 32'h0 : _GEN_5148;
  assign _GEN_5150 = 9'h55 == _T_82861 ? 32'h0 : _GEN_5149;
  assign _GEN_5151 = 9'h56 == _T_82861 ? 32'h0 : _GEN_5150;
  assign _GEN_5152 = 9'h57 == _T_82861 ? 32'h0 : _GEN_5151;
  assign _GEN_5153 = 9'h58 == _T_82861 ? 32'h0 : _GEN_5152;
  assign _GEN_5154 = 9'h59 == _T_82861 ? 32'h0 : _GEN_5153;
  assign _GEN_5155 = 9'h5a == _T_82861 ? 32'h0 : _GEN_5154;
  assign _GEN_5156 = 9'h5b == _T_82861 ? 32'h0 : _GEN_5155;
  assign _GEN_5157 = 9'h5c == _T_82861 ? 32'h0 : _GEN_5156;
  assign _GEN_5158 = 9'h5d == _T_82861 ? 32'h0 : _GEN_5157;
  assign _GEN_5159 = 9'h5e == _T_82861 ? 32'h0 : _GEN_5158;
  assign _GEN_5160 = 9'h5f == _T_82861 ? 32'h0 : _GEN_5159;
  assign _GEN_5161 = 9'h60 == _T_82861 ? 32'h0 : _GEN_5160;
  assign _GEN_5162 = 9'h61 == _T_82861 ? 32'h0 : _GEN_5161;
  assign _GEN_5163 = 9'h62 == _T_82861 ? 32'h0 : _GEN_5162;
  assign _GEN_5164 = 9'h63 == _T_82861 ? 32'h0 : _GEN_5163;
  assign _GEN_5165 = 9'h64 == _T_82861 ? 32'h0 : _GEN_5164;
  assign _GEN_5166 = 9'h65 == _T_82861 ? 32'h0 : _GEN_5165;
  assign _GEN_5167 = 9'h66 == _T_82861 ? 32'h0 : _GEN_5166;
  assign _GEN_5168 = 9'h67 == _T_82861 ? 32'h0 : _GEN_5167;
  assign _GEN_5169 = 9'h68 == _T_82861 ? 32'h0 : _GEN_5168;
  assign _GEN_5170 = 9'h69 == _T_82861 ? 32'h0 : _GEN_5169;
  assign _GEN_5171 = 9'h6a == _T_82861 ? 32'h0 : _GEN_5170;
  assign _GEN_5172 = 9'h6b == _T_82861 ? 32'h0 : _GEN_5171;
  assign _GEN_5173 = 9'h6c == _T_82861 ? 32'h0 : _GEN_5172;
  assign _GEN_5174 = 9'h6d == _T_82861 ? 32'h0 : _GEN_5173;
  assign _GEN_5175 = 9'h6e == _T_82861 ? 32'h0 : _GEN_5174;
  assign _GEN_5176 = 9'h6f == _T_82861 ? 32'h0 : _GEN_5175;
  assign _GEN_5177 = 9'h70 == _T_82861 ? 32'h0 : _GEN_5176;
  assign _GEN_5178 = 9'h71 == _T_82861 ? 32'h0 : _GEN_5177;
  assign _GEN_5179 = 9'h72 == _T_82861 ? 32'h0 : _GEN_5178;
  assign _GEN_5180 = 9'h73 == _T_82861 ? 32'h0 : _GEN_5179;
  assign _GEN_5181 = 9'h74 == _T_82861 ? 32'h0 : _GEN_5180;
  assign _GEN_5182 = 9'h75 == _T_82861 ? 32'h0 : _GEN_5181;
  assign _GEN_5183 = 9'h76 == _T_82861 ? 32'h0 : _GEN_5182;
  assign _GEN_5184 = 9'h77 == _T_82861 ? 32'h0 : _GEN_5183;
  assign _GEN_5185 = 9'h78 == _T_82861 ? 32'h0 : _GEN_5184;
  assign _GEN_5186 = 9'h79 == _T_82861 ? 32'h0 : _GEN_5185;
  assign _GEN_5187 = 9'h7a == _T_82861 ? 32'h0 : _GEN_5186;
  assign _GEN_5188 = 9'h7b == _T_82861 ? 32'h0 : _GEN_5187;
  assign _GEN_5189 = 9'h7c == _T_82861 ? 32'h0 : _GEN_5188;
  assign _GEN_5190 = 9'h7d == _T_82861 ? 32'h0 : _GEN_5189;
  assign _GEN_5191 = 9'h7e == _T_82861 ? 32'h0 : _GEN_5190;
  assign _GEN_5192 = 9'h7f == _T_82861 ? 32'h0 : _GEN_5191;
  assign _GEN_5193 = 9'h80 == _T_82861 ? 32'h0 : _GEN_5192;
  assign _GEN_5194 = 9'h81 == _T_82861 ? 32'h0 : _GEN_5193;
  assign _GEN_5195 = 9'h82 == _T_82861 ? 32'h0 : _GEN_5194;
  assign _GEN_5196 = 9'h83 == _T_82861 ? 32'h0 : _GEN_5195;
  assign _GEN_5197 = 9'h84 == _T_82861 ? 32'h0 : _GEN_5196;
  assign _GEN_5198 = 9'h85 == _T_82861 ? 32'h0 : _GEN_5197;
  assign _GEN_5199 = 9'h86 == _T_82861 ? 32'h0 : _GEN_5198;
  assign _GEN_5200 = 9'h87 == _T_82861 ? 32'h0 : _GEN_5199;
  assign _GEN_5201 = 9'h88 == _T_82861 ? 32'h0 : _GEN_5200;
  assign _GEN_5202 = 9'h89 == _T_82861 ? 32'h0 : _GEN_5201;
  assign _GEN_5203 = 9'h8a == _T_82861 ? 32'h0 : _GEN_5202;
  assign _GEN_5204 = 9'h8b == _T_82861 ? 32'h0 : _GEN_5203;
  assign _GEN_5205 = 9'h8c == _T_82861 ? 32'h0 : _GEN_5204;
  assign _GEN_5206 = 9'h8d == _T_82861 ? 32'h0 : _GEN_5205;
  assign _GEN_5207 = 9'h8e == _T_82861 ? 32'h0 : _GEN_5206;
  assign _GEN_5208 = 9'h8f == _T_82861 ? 32'h0 : _GEN_5207;
  assign _GEN_5209 = 9'h90 == _T_82861 ? 32'h0 : _GEN_5208;
  assign _GEN_5210 = 9'h91 == _T_82861 ? 32'h0 : _GEN_5209;
  assign _GEN_5211 = 9'h92 == _T_82861 ? 32'h0 : _GEN_5210;
  assign _GEN_5212 = 9'h93 == _T_82861 ? 32'h0 : _GEN_5211;
  assign _GEN_5213 = 9'h94 == _T_82861 ? 32'h0 : _GEN_5212;
  assign _GEN_5214 = 9'h95 == _T_82861 ? 32'h0 : _GEN_5213;
  assign _GEN_5215 = 9'h96 == _T_82861 ? 32'h0 : _GEN_5214;
  assign _GEN_5216 = 9'h97 == _T_82861 ? 32'h0 : _GEN_5215;
  assign _GEN_5217 = 9'h98 == _T_82861 ? 32'h0 : _GEN_5216;
  assign _GEN_5218 = 9'h99 == _T_82861 ? 32'h0 : _GEN_5217;
  assign _GEN_5219 = 9'h9a == _T_82861 ? 32'h0 : _GEN_5218;
  assign _GEN_5220 = 9'h9b == _T_82861 ? 32'h0 : _GEN_5219;
  assign _GEN_5221 = 9'h9c == _T_82861 ? 32'h0 : _GEN_5220;
  assign _GEN_5222 = 9'h9d == _T_82861 ? 32'h0 : _GEN_5221;
  assign _GEN_5223 = 9'h9e == _T_82861 ? 32'h0 : _GEN_5222;
  assign _GEN_5224 = 9'h9f == _T_82861 ? 32'h0 : _GEN_5223;
  assign _GEN_5225 = 9'ha0 == _T_82861 ? 32'h0 : _GEN_5224;
  assign _GEN_5226 = 9'ha1 == _T_82861 ? 32'h0 : _GEN_5225;
  assign _GEN_5227 = 9'ha2 == _T_82861 ? 32'h0 : _GEN_5226;
  assign _GEN_5228 = 9'ha3 == _T_82861 ? 32'h0 : _GEN_5227;
  assign _GEN_5229 = 9'ha4 == _T_82861 ? 32'h0 : _GEN_5228;
  assign _GEN_5230 = 9'ha5 == _T_82861 ? 32'h0 : _GEN_5229;
  assign _GEN_5231 = 9'ha6 == _T_82861 ? 32'h0 : _GEN_5230;
  assign _GEN_5232 = 9'ha7 == _T_82861 ? 32'h0 : _GEN_5231;
  assign _GEN_5233 = 9'ha8 == _T_82861 ? 32'h0 : _GEN_5232;
  assign _GEN_5234 = 9'ha9 == _T_82861 ? 32'h0 : _GEN_5233;
  assign _GEN_5235 = 9'haa == _T_82861 ? 32'h0 : _GEN_5234;
  assign _GEN_5236 = 9'hab == _T_82861 ? 32'h0 : _GEN_5235;
  assign _GEN_5237 = 9'hac == _T_82861 ? 32'h0 : _GEN_5236;
  assign _GEN_5238 = 9'had == _T_82861 ? 32'h0 : _GEN_5237;
  assign _GEN_5239 = 9'hae == _T_82861 ? 32'h0 : _GEN_5238;
  assign _GEN_5240 = 9'haf == _T_82861 ? 32'h0 : _GEN_5239;
  assign _GEN_5241 = 9'hb0 == _T_82861 ? 32'h0 : _GEN_5240;
  assign _GEN_5242 = 9'hb1 == _T_82861 ? 32'h0 : _GEN_5241;
  assign _GEN_5243 = 9'hb2 == _T_82861 ? 32'h0 : _GEN_5242;
  assign _GEN_5244 = 9'hb3 == _T_82861 ? 32'h0 : _GEN_5243;
  assign _GEN_5245 = 9'hb4 == _T_82861 ? 32'h0 : _GEN_5244;
  assign _GEN_5246 = 9'hb5 == _T_82861 ? 32'h0 : _GEN_5245;
  assign _GEN_5247 = 9'hb6 == _T_82861 ? 32'h0 : _GEN_5246;
  assign _GEN_5248 = 9'hb7 == _T_82861 ? 32'h0 : _GEN_5247;
  assign _GEN_5249 = 9'hb8 == _T_82861 ? 32'h0 : _GEN_5248;
  assign _GEN_5250 = 9'hb9 == _T_82861 ? 32'h0 : _GEN_5249;
  assign _GEN_5251 = 9'hba == _T_82861 ? 32'h0 : _GEN_5250;
  assign _GEN_5252 = 9'hbb == _T_82861 ? 32'h0 : _GEN_5251;
  assign _GEN_5253 = 9'hbc == _T_82861 ? 32'h0 : _GEN_5252;
  assign _GEN_5254 = 9'hbd == _T_82861 ? 32'h0 : _GEN_5253;
  assign _GEN_5255 = 9'hbe == _T_82861 ? 32'h0 : _GEN_5254;
  assign _GEN_5256 = 9'hbf == _T_82861 ? 32'h0 : _GEN_5255;
  assign _GEN_5257 = 9'hc0 == _T_82861 ? 32'h380006f : _GEN_5256;
  assign _GEN_5258 = 9'hc1 == _T_82861 ? 32'h0 : _GEN_5257;
  assign _GEN_5259 = 9'hc2 == _T_82861 ? 32'h0 : _GEN_5258;
  assign _GEN_5260 = 9'hc3 == _T_82861 ? 32'h0 : _GEN_5259;
  assign _GEN_5261 = 9'hc4 == _T_82861 ? 32'h0 : _GEN_5260;
  assign _GEN_5262 = 9'hc5 == _T_82861 ? 32'h0 : _GEN_5261;
  assign _GEN_5263 = 9'hc6 == _T_82861 ? 32'h0 : _GEN_5262;
  assign _GEN_5264 = 9'hc7 == _T_82861 ? 32'h0 : _GEN_5263;
  assign _GEN_5265 = 9'hc8 == _T_82861 ? 32'h0 : _GEN_5264;
  assign _GEN_5266 = 9'hc9 == _T_82861 ? 32'h0 : _GEN_5265;
  assign _GEN_5267 = 9'hca == _T_82861 ? 32'h0 : _GEN_5266;
  assign _GEN_5268 = 9'hcb == _T_82861 ? 32'h0 : _GEN_5267;
  assign _GEN_5269 = 9'hcc == _T_82861 ? 32'h0 : _GEN_5268;
  assign _GEN_5270 = 9'hcd == _T_82861 ? 32'h0 : _GEN_5269;
  assign _GEN_5271 = 9'hce == _T_82861 ? abstractGeneratedMem_0 : _GEN_5270;
  assign _GEN_5272 = 9'hcf == _T_82861 ? abstractGeneratedMem_1 : _GEN_5271;
  assign _GEN_5273 = 9'hd0 == _T_82861 ? _T_4738 : _GEN_5272;
  assign _GEN_5274 = 9'hd1 == _T_82861 ? _T_4418 : _GEN_5273;
  assign _GEN_5275 = 9'hd2 == _T_82861 ? _T_4898 : _GEN_5274;
  assign _GEN_5276 = 9'hd3 == _T_82861 ? _T_5658 : _GEN_5275;
  assign _GEN_5277 = 9'hd4 == _T_82861 ? _T_6218 : _GEN_5276;
  assign _GEN_5278 = 9'hd5 == _T_82861 ? _T_3938 : _GEN_5277;
  assign _GEN_5279 = 9'hd6 == _T_82861 ? _T_4258 : _GEN_5278;
  assign _GEN_5280 = 9'hd7 == _T_82861 ? _T_5498 : _GEN_5279;
  assign _GEN_5281 = 9'hd8 == _T_82861 ? _T_6018 : _GEN_5280;
  assign _GEN_5282 = 9'hd9 == _T_82861 ? _T_4578 : _GEN_5281;
  assign _GEN_5283 = 9'hda == _T_82861 ? _T_3738 : _GEN_5282;
  assign _GEN_5284 = 9'hdb == _T_82861 ? _T_5858 : _GEN_5283;
  assign _GEN_5285 = 9'hdc == _T_82861 ? _T_5338 : _GEN_5284;
  assign _GEN_5286 = 9'hdd == _T_82861 ? _T_5058 : _GEN_5285;
  assign _GEN_5287 = 9'hde == _T_82861 ? _T_4098 : _GEN_5286;
  assign _GEN_5288 = 9'hdf == _T_82861 ? _T_6578 : _GEN_5287;
  assign _GEN_5289 = 9'he0 == _T_82861 ? _T_6418 : _GEN_5288;
  assign _GEN_5290 = 9'he1 == _T_82861 ? 32'h0 : _GEN_5289;
  assign _GEN_5291 = 9'he2 == _T_82861 ? 32'h0 : _GEN_5290;
  assign _GEN_5292 = 9'he3 == _T_82861 ? 32'h0 : _GEN_5291;
  assign _GEN_5293 = 9'he4 == _T_82861 ? 32'h0 : _GEN_5292;
  assign _GEN_5294 = 9'he5 == _T_82861 ? 32'h0 : _GEN_5293;
  assign _GEN_5295 = 9'he6 == _T_82861 ? 32'h0 : _GEN_5294;
  assign _GEN_5296 = 9'he7 == _T_82861 ? 32'h0 : _GEN_5295;
  assign _GEN_5297 = 9'he8 == _T_82861 ? 32'h0 : _GEN_5296;
  assign _GEN_5298 = 9'he9 == _T_82861 ? 32'h0 : _GEN_5297;
  assign _GEN_5299 = 9'hea == _T_82861 ? 32'h0 : _GEN_5298;
  assign _GEN_5300 = 9'heb == _T_82861 ? 32'h0 : _GEN_5299;
  assign _GEN_5301 = 9'hec == _T_82861 ? 32'h0 : _GEN_5300;
  assign _GEN_5302 = 9'hed == _T_82861 ? 32'h0 : _GEN_5301;
  assign _GEN_5303 = 9'hee == _T_82861 ? 32'h0 : _GEN_5302;
  assign _GEN_5304 = 9'hef == _T_82861 ? 32'h0 : _GEN_5303;
  assign _GEN_5305 = 9'hf0 == _T_82861 ? 32'h0 : _GEN_5304;
  assign _GEN_5306 = 9'hf1 == _T_82861 ? 32'h0 : _GEN_5305;
  assign _GEN_5307 = 9'hf2 == _T_82861 ? 32'h0 : _GEN_5306;
  assign _GEN_5308 = 9'hf3 == _T_82861 ? 32'h0 : _GEN_5307;
  assign _GEN_5309 = 9'hf4 == _T_82861 ? 32'h0 : _GEN_5308;
  assign _GEN_5310 = 9'hf5 == _T_82861 ? 32'h0 : _GEN_5309;
  assign _GEN_5311 = 9'hf6 == _T_82861 ? 32'h0 : _GEN_5310;
  assign _GEN_5312 = 9'hf7 == _T_82861 ? 32'h0 : _GEN_5311;
  assign _GEN_5313 = 9'hf8 == _T_82861 ? 32'h0 : _GEN_5312;
  assign _GEN_5314 = 9'hf9 == _T_82861 ? 32'h0 : _GEN_5313;
  assign _GEN_5315 = 9'hfa == _T_82861 ? 32'h0 : _GEN_5314;
  assign _GEN_5316 = 9'hfb == _T_82861 ? 32'h0 : _GEN_5315;
  assign _GEN_5317 = 9'hfc == _T_82861 ? 32'h0 : _GEN_5316;
  assign _GEN_5318 = 9'hfd == _T_82861 ? 32'h0 : _GEN_5317;
  assign _GEN_5319 = 9'hfe == _T_82861 ? 32'h0 : _GEN_5318;
  assign _GEN_5320 = 9'hff == _T_82861 ? 32'h0 : _GEN_5319;
  assign _GEN_5321 = 9'h100 == _T_82861 ? _T_53243 : _GEN_5320;
  assign _GEN_5322 = 9'h101 == _T_82861 ? _T_40003 : _GEN_5321;
  assign _GEN_5323 = 9'h102 == _T_82861 ? _T_73203 : _GEN_5322;
  assign _GEN_5324 = 9'h103 == _T_82861 ? _T_58723 : _GEN_5323;
  assign _GEN_5325 = 9'h104 == _T_82861 ? _T_48523 : _GEN_5324;
  assign _GEN_5326 = 9'h105 == _T_82861 ? _T_42243 : _GEN_5325;
  assign _GEN_5327 = 9'h106 == _T_82861 ? _T_76443 : _GEN_5326;
  assign _GEN_5328 = 9'h107 == _T_82861 ? _T_69003 : _GEN_5327;
  assign _GEN_5329 = 9'h108 == _T_82861 ? _T_57083 : _GEN_5328;
  assign _GEN_5330 = 9'h109 == _T_82861 ? _T_45603 : _GEN_5329;
  assign _GEN_5331 = 9'h10a == _T_82861 ? _T_55323 : _GEN_5330;
  assign _GEN_5332 = 9'h10b == _T_82861 ? _T_65643 : _GEN_5331;
  assign _GEN_5333 = 9'h10c == _T_82861 ? _T_78203 : _GEN_5332;
  assign _GEN_5334 = 9'h10d == _T_82861 ? _T_37923 : _GEN_5333;
  assign _GEN_5335 = 9'h10e == _T_82861 ? _T_47243 : _GEN_5334;
  assign _GEN_5336 = 9'h10f == _T_82861 ? _T_62083 : _GEN_5335;
  assign _GEN_5337 = 9'h110 == _T_82861 ? _T_74843 : _GEN_5336;
  assign _GEN_5338 = 9'h111 == _T_82861 ? _T_76923 : _GEN_5337;
  assign _GEN_5339 = 9'h112 == _T_82861 ? _T_60643 : _GEN_5338;
  assign _GEN_5340 = 9'h113 == _T_82861 ? _T_49683 : _GEN_5339;
  assign _GEN_5341 = 9'h114 == _T_82861 ? _T_36963 : _GEN_5340;
  assign _GEN_5342 = 9'h115 == _T_82861 ? _T_80443 : _GEN_5341;
  assign _GEN_5343 = 9'h116 == _T_82861 ? _T_64683 : _GEN_5342;
  assign _GEN_5344 = 9'h117 == _T_82861 ? _T_57243 : _GEN_5343;
  assign _GEN_5345 = 9'h118 == _T_82861 ? _T_44483 : _GEN_5344;
  assign _GEN_5346 = 9'h119 == _T_82861 ? _T_58563 : _GEN_5345;
  assign _GEN_5347 = 9'h11a == _T_82861 ? _T_68363 : _GEN_5346;
  assign _GEN_5348 = 9'h11b == _T_82861 ? _T_79163 : _GEN_5347;
  assign _GEN_5349 = 9'h11c == _T_82861 ? _T_41283 : _GEN_5348;
  assign _GEN_5350 = 9'h11d == _T_82861 ? _T_51483 : _GEN_5349;
  assign _GEN_5351 = 9'h11e == _T_82861 ? _T_58243 : _GEN_5350;
  assign _GEN_5352 = 9'h11f == _T_82861 ? _T_75483 : _GEN_5351;
  assign _GEN_5353 = 9'h120 == _T_82861 ? _T_39363 : _GEN_5352;
  assign _GEN_5354 = 9'h121 == _T_82861 ? _T_41763 : _GEN_5353;
  assign _GEN_5355 = 9'h122 == _T_82861 ? _T_74003 : _GEN_5354;
  assign _GEN_5356 = 9'h123 == _T_82861 ? _T_58403 : _GEN_5355;
  assign _GEN_5357 = 9'h124 == _T_82861 ? _T_46443 : _GEN_5356;
  assign _GEN_5358 = 9'h125 == _T_82861 ? _T_44803 : _GEN_5357;
  assign _GEN_5359 = 9'h126 == _T_82861 ? _T_77723 : _GEN_5358;
  assign _GEN_5360 = 9'h127 == _T_82861 ? _T_68203 : _GEN_5359;
  assign _GEN_5361 = 9'h128 == _T_82861 ? _T_57443 : _GEN_5360;
  assign _GEN_5362 = 9'h129 == _T_82861 ? _T_49003 : _GEN_5361;
  assign _GEN_5363 = 9'h12a == _T_82861 ? _T_56283 : _GEN_5362;
  assign _GEN_5364 = 9'h12b == _T_82861 ? _T_65483 : _GEN_5363;
  assign _GEN_5365 = 9'h12c == _T_82861 ? _T_75643 : _GEN_5364;
  assign _GEN_5366 = 9'h12d == _T_82861 ? _T_39523 : _GEN_5365;
  assign _GEN_5367 = 9'h12e == _T_82861 ? _T_48363 : _GEN_5366;
  assign _GEN_5368 = 9'h12f == _T_82861 ? _T_61923 : _GEN_5367;
  assign _GEN_5369 = 9'h130 == _T_82861 ? _T_73043 : _GEN_5368;
  assign _GEN_5370 = 9'h131 == _T_82861 ? _T_77243 : _GEN_5369;
  assign _GEN_5371 = 9'h132 == _T_82861 ? _T_65323 : _GEN_5370;
  assign _GEN_5372 = 9'h133 == _T_82861 ? _T_46283 : _GEN_5371;
  assign _GEN_5373 = 9'h134 == _T_82861 ? _T_37123 : _GEN_5372;
  assign _GEN_5374 = 9'h135 == _T_82861 ? _T_81883 : _GEN_5373;
  assign _GEN_5375 = 9'h136 == _T_82861 ? _T_69163 : _GEN_5374;
  assign _GEN_5376 = 9'h137 == _T_82861 ? _T_55803 : _GEN_5375;
  assign _GEN_5377 = 9'h138 == _T_82861 ? _T_46083 : _GEN_5376;
  assign _GEN_5378 = 9'h139 == _T_82861 ? _T_59523 : _GEN_5377;
  assign _GEN_5379 = 9'h13a == _T_82861 ? _T_70963 : _GEN_5378;
  assign _GEN_5380 = 9'h13b == _T_82861 ? _T_75963 : _GEN_5379;
  assign _GEN_5381 = 9'h13c == _T_82861 ? _T_42083 : _GEN_5380;
  assign _GEN_5382 = 9'h13d == _T_82861 ? _T_51963 : _GEN_5381;
  assign _GEN_5383 = 9'h13e == _T_82861 ? _T_61443 : _GEN_5382;
  assign _GEN_5384 = 9'h13f == _T_82861 ? _T_72883 : _GEN_5383;
  assign _GEN_5385 = 9'h140 == _T_82861 ? _T_39683 : _GEN_5384;
  assign _GEN_5386 = 9'h141 == _T_82861 ? _T_43043 : _GEN_5385;
  assign _GEN_5387 = 9'h142 == _T_82861 ? _T_81083 : _GEN_5386;
  assign _GEN_5388 = 9'h143 == _T_82861 ? _T_63363 : _GEN_5387;
  assign _GEN_5389 = 9'h144 == _T_82861 ? _T_51323 : _GEN_5388;
  assign _GEN_5390 = 9'h145 == _T_82861 ? _T_41603 : _GEN_5389;
  assign _GEN_5391 = 9'h146 == _T_82861 ? _T_77563 : _GEN_5390;
  assign _GEN_5392 = 9'h147 == _T_82861 ? _T_68683 : _GEN_5391;
  assign _GEN_5393 = 9'h148 == _T_82861 ? _T_52923 : _GEN_5392;
  assign _GEN_5394 = 9'h149 == _T_82861 ? _T_50523 : _GEN_5393;
  assign _GEN_5395 = 9'h14a == _T_82861 ? _T_64043 : _GEN_5394;
  assign _GEN_5396 = 9'h14b == _T_82861 ? _T_69363 : _GEN_5395;
  assign _GEN_5397 = 9'h14c == _T_82861 ? _T_79803 : _GEN_5396;
  assign _GEN_5398 = 9'h14d == _T_82861 ? _T_35683 : _GEN_5397;
  assign _GEN_5399 = 9'h14e == _T_82861 ? _T_48203 : _GEN_5398;
  assign _GEN_5400 = 9'h14f == _T_82861 ? _T_60003 : _GEN_5399;
  assign _GEN_5401 = 9'h150 == _T_82861 ? _T_70643 : _GEN_5400;
  assign _GEN_5402 = 9'h151 == _T_82861 ? _T_81403 : _GEN_5401;
  assign _GEN_5403 = 9'h152 == _T_82861 ? _T_70163 : _GEN_5402;
  assign _GEN_5404 = 9'h153 == _T_82861 ? _T_53563 : _GEN_5403;
  assign _GEN_5405 = 9'h154 == _T_82861 ? _T_38883 : _GEN_5404;
  assign _GEN_5406 = 9'h155 == _T_82861 ? _T_77883 : _GEN_5405;
  assign _GEN_5407 = 9'h156 == _T_82861 ? _T_67563 : _GEN_5406;
  assign _GEN_5408 = 9'h157 == _T_82861 ? _T_55163 : _GEN_5407;
  assign _GEN_5409 = 9'h158 == _T_82861 ? _T_40643 : _GEN_5408;
  assign _GEN_5410 = 9'h159 == _T_82861 ? _T_62883 : _GEN_5409;
  assign _GEN_5411 = 9'h15a == _T_82861 ? _T_75163 : _GEN_5410;
  assign _GEN_5412 = 9'h15b == _T_82861 ? _T_35523 : _GEN_5411;
  assign _GEN_5413 = 9'h15c == _T_82861 ? _T_43843 : _GEN_5412;
  assign _GEN_5414 = 9'h15d == _T_82861 ? _T_48683 : _GEN_5413;
  assign _GEN_5415 = 9'h15e == _T_82861 ? _T_60163 : _GEN_5414;
  assign _GEN_5416 = 9'h15f == _T_82861 ? _T_73363 : _GEN_5415;
  assign _GEN_5417 = 9'h160 == _T_82861 ? _T_36323 : _GEN_5416;
  assign _GEN_5418 = 9'h161 == _T_82861 ? _T_44003 : _GEN_5417;
  assign _GEN_5419 = 9'h162 == _T_82861 ? _T_81723 : _GEN_5418;
  assign _GEN_5420 = 9'h163 == _T_82861 ? _T_67723 : _GEN_5419;
  assign _GEN_5421 = 9'h164 == _T_82861 ? _T_52443 : _GEN_5420;
  assign _GEN_5422 = 9'h165 == _T_82861 ? _T_40803 : _GEN_5421;
  assign _GEN_5423 = 9'h166 == _T_82861 ? _T_78363 : _GEN_5422;
  assign _GEN_5424 = 9'h167 == _T_82861 ? _T_70483 : _GEN_5423;
  assign _GEN_5425 = 9'h168 == _T_82861 ? _T_55483 : _GEN_5424;
  assign _GEN_5426 = 9'h169 == _T_82861 ? _T_50163 : _GEN_5425;
  assign _GEN_5427 = 9'h16a == _T_82861 ? _T_61123 : _GEN_5426;
  assign _GEN_5428 = 9'h16b == _T_82861 ? _T_71763 : _GEN_5427;
  assign _GEN_5429 = 9'h16c == _T_82861 ? _T_82843 : _GEN_5428;
  assign _GEN_5430 = 9'h16d == _T_82861 ? _T_35203 : _GEN_5429;
  assign _GEN_5431 = 9'h16e == _T_82861 ? _T_47883 : _GEN_5430;
  assign _GEN_5432 = 9'h16f == _T_82861 ? _T_63043 : _GEN_5431;
  assign _GEN_5433 = 9'h170 == _T_82861 ? _T_72563 : _GEN_5432;
  assign _GEN_5434 = 9'h171 == _T_82861 ? _T_80923 : _GEN_5433;
  assign _GEN_5435 = 9'h172 == _T_82861 ? _T_69683 : _GEN_5434;
  assign _GEN_5436 = 9'h173 == _T_82861 ? _T_54843 : _GEN_5435;
  assign _GEN_5437 = 9'h174 == _T_82861 ? _T_40323 : _GEN_5436;
  assign _GEN_5438 = 9'h175 == _T_82861 ? _T_77083 : _GEN_5437;
  assign _GEN_5439 = 9'h176 == _T_82861 ? _T_66923 : _GEN_5438;
  assign _GEN_5440 = 9'h177 == _T_82861 ? _T_57763 : _GEN_5439;
  assign _GEN_5441 = 9'h178 == _T_82861 ? _T_43203 : _GEN_5440;
  assign _GEN_5442 = 9'h179 == _T_82861 ? _T_60963 : _GEN_5441;
  assign _GEN_5443 = 9'h17a == _T_82861 ? _T_74163 : _GEN_5442;
  assign _GEN_5444 = 9'h17b == _T_82861 ? _T_37443 : _GEN_5443;
  assign _GEN_5445 = 9'h17c == _T_82861 ? _T_46763 : _GEN_5444;
  assign _GEN_5446 = 9'h17d == _T_82861 ? _T_47563 : _GEN_5445;
  assign _GEN_5447 = 9'h17e == _T_82861 ? _T_59363 : _GEN_5446;
  assign _GEN_5448 = 9'h17f == _T_82861 ? _T_75003 : _GEN_5447;
  assign _GEN_5449 = 9'h180 == _T_82861 ? _T_38243 : _GEN_5448;
  assign _GEN_5450 = 9'h181 == _T_82861 ? _T_38083 : _GEN_5449;
  assign _GEN_5451 = 9'h182 == _T_82861 ? _T_70803 : _GEN_5450;
  assign _GEN_5452 = 9'h183 == _T_82861 ? _T_62563 : _GEN_5451;
  assign _GEN_5453 = 9'h184 == _T_82861 ? _T_52283 : _GEN_5452;
  assign _GEN_5454 = 9'h185 == _T_82861 ? _T_40163 : _GEN_5453;
  assign _GEN_5455 = 9'h186 == _T_82861 ? _T_73523 : _GEN_5454;
  assign _GEN_5456 = 9'h187 == _T_82861 ? _T_59043 : _GEN_5455;
  assign _GEN_5457 = 9'h188 == _T_82861 ? _T_48843 : _GEN_5456;
  assign _GEN_5458 = 9'h189 == _T_82861 ? _T_54363 : _GEN_5457;
  assign _GEN_5459 = 9'h18a == _T_82861 ? _T_65163 : _GEN_5458;
  assign _GEN_5460 = 9'h18b == _T_82861 ? _T_79483 : _GEN_5459;
  assign _GEN_5461 = 9'h18c == _T_82861 ? _T_45123 : _GEN_5460;
  assign _GEN_5462 = 9'h18d == _T_82861 ? _T_44323 : _GEN_5461;
  assign _GEN_5463 = 9'h18e == _T_82861 ? _T_55963 : _GEN_5462;
  assign _GEN_5464 = 9'h18f == _T_82861 ? _T_64523 : _GEN_5463;
  assign _GEN_5465 = 9'h190 == _T_82861 ? _T_78843 : _GEN_5464;
  assign _GEN_5466 = 9'h191 == _T_82861 ? _T_73683 : _GEN_5465;
  assign _GEN_5467 = 9'h192 == _T_82861 ? _T_58083 : _GEN_5466;
  assign _GEN_5468 = 9'h193 == _T_82861 ? _T_52123 : _GEN_5467;
  assign _GEN_5469 = 9'h194 == _T_82861 ? _T_39043 : _GEN_5468;
  assign _GEN_5470 = 9'h195 == _T_82861 ? _T_76603 : _GEN_5469;
  assign _GEN_5471 = 9'h196 == _T_82861 ? _T_60323 : _GEN_5470;
  assign _GEN_5472 = 9'h197 == _T_82861 ? _T_49363 : _GEN_5471;
  assign _GEN_5473 = 9'h198 == _T_82861 ? _T_36483 : _GEN_5472;
  assign _GEN_5474 = 9'h199 == _T_82861 ? _T_68843 : _GEN_5473;
  assign _GEN_5475 = 9'h19a == _T_82861 ? _T_76283 : _GEN_5474;
  assign _GEN_5476 = 9'h19b == _T_82861 ? _T_45283 : _GEN_5475;
  assign _GEN_5477 = 9'h19c == _T_82861 ? _T_56443 : _GEN_5476;
  assign _GEN_5478 = 9'h19d == _T_82861 ? _T_58883 : _GEN_5477;
  assign _GEN_5479 = 9'h19e == _T_82861 ? _T_68523 : _GEN_5478;
  assign _GEN_5480 = 9'h19f == _T_82861 ? _T_79323 : _GEN_5479;
  assign _GEN_5481 = 9'h1a0 == _T_82861 ? _T_41443 : _GEN_5480;
  assign _GEN_5482 = 9'h1a1 == _T_82861 ? _T_39203 : _GEN_5481;
  assign _GEN_5483 = 9'h1a2 == _T_82861 ? _T_73843 : _GEN_5482;
  assign _GEN_5484 = 9'h1a3 == _T_82861 ? _T_60803 : _GEN_5483;
  assign _GEN_5485 = 9'h1a4 == _T_82861 ? _T_52603 : _GEN_5484;
  assign _GEN_5486 = 9'h1a5 == _T_82861 ? _T_41123 : _GEN_5485;
  assign _GEN_5487 = 9'h1a6 == _T_82861 ? _T_76763 : _GEN_5486;
  assign _GEN_5488 = 9'h1a7 == _T_82861 ? _T_57923 : _GEN_5487;
  assign _GEN_5489 = 9'h1a8 == _T_82861 ? _T_49163 : _GEN_5488;
  assign _GEN_5490 = 9'h1a9 == _T_82861 ? _T_56603 : _GEN_5489;
  assign _GEN_5491 = 9'h1aa == _T_82861 ? _T_66603 : _GEN_5490;
  assign _GEN_5492 = 9'h1ab == _T_82861 ? _T_79963 : _GEN_5491;
  assign _GEN_5493 = 9'h1ac == _T_82861 ? _T_45443 : _GEN_5492;
  assign _GEN_5494 = 9'h1ad == _T_82861 ? _T_49523 : _GEN_5493;
  assign _GEN_5495 = 9'h1ae == _T_82861 ? _T_56923 : _GEN_5494;
  assign _GEN_5496 = 9'h1af == _T_82861 ? _T_66123 : _GEN_5495;
  assign _GEN_5497 = 9'h1b0 == _T_82861 ? _T_76123 : _GEN_5496;
  assign _GEN_5498 = 9'h1b1 == _T_82861 ? _T_74323 : _GEN_5497;
  assign _GEN_5499 = 9'h1b2 == _T_82861 ? _T_61763 : _GEN_5498;
  assign _GEN_5500 = 9'h1b3 == _T_82861 ? _T_50363 : _GEN_5499;
  assign _GEN_5501 = 9'h1b4 == _T_82861 ? _T_39843 : _GEN_5500;
  assign _GEN_5502 = 9'h1b5 == _T_82861 ? _T_78523 : _GEN_5501;
  assign _GEN_5503 = 9'h1b6 == _T_82861 ? _T_65963 : _GEN_5502;
  assign _GEN_5504 = 9'h1b7 == _T_82861 ? _T_47083 : _GEN_5503;
  assign _GEN_5505 = 9'h1b8 == _T_82861 ? _T_37603 : _GEN_5504;
  assign _GEN_5506 = 9'h1b9 == _T_82861 ? _T_69523 : _GEN_5505;
  assign _GEN_5507 = 9'h1ba == _T_82861 ? _T_80603 : _GEN_5506;
  assign _GEN_5508 = 9'h1bb == _T_82861 ? _T_42883 : _GEN_5507;
  assign _GEN_5509 = 9'h1bc == _T_82861 ? _T_57603 : _GEN_5508;
  assign _GEN_5510 = 9'h1bd == _T_82861 ? _T_59203 : _GEN_5509;
  assign _GEN_5511 = 9'h1be == _T_82861 ? _T_71123 : _GEN_5510;
  assign _GEN_5512 = 9'h1bf == _T_82861 ? _T_75803 : _GEN_5511;
  assign _GEN_5513 = 9'h1c0 == _T_82861 ? _T_41923 : _GEN_5512;
  assign _GEN_5514 = 9'h1c1 == _T_82861 ? _T_37283 : _GEN_5513;
  assign _GEN_5515 = 9'h1c2 == _T_82861 ? _T_71603 : _GEN_5514;
  assign _GEN_5516 = 9'h1c3 == _T_82861 ? _T_61283 : _GEN_5515;
  assign _GEN_5517 = 9'h1c4 == _T_82861 ? _T_46603 : _GEN_5516;
  assign _GEN_5518 = 9'h1c5 == _T_82861 ? _T_44963 : _GEN_5517;
  assign _GEN_5519 = 9'h1c6 == _T_82861 ? _T_82683 : _GEN_5518;
  assign _GEN_5520 = 9'h1c7 == _T_82861 ? _T_64843 : _GEN_5519;
  assign _GEN_5521 = 9'h1c8 == _T_82861 ? _T_51163 : _GEN_5520;
  assign _GEN_5522 = 9'h1c9 == _T_82861 ? _T_54683 : _GEN_5521;
  assign _GEN_5523 = 9'h1ca == _T_82861 ? _T_67883 : _GEN_5522;
  assign _GEN_5524 = 9'h1cb == _T_82861 ? _T_80283 : _GEN_5523;
  assign _GEN_5525 = 9'h1cc == _T_82861 ? _T_40963 : _GEN_5524;
  assign _GEN_5526 = 9'h1cd == _T_82861 ? _T_50843 : _GEN_5525;
  assign _GEN_5527 = 9'h1ce == _T_82861 ? _T_64203 : _GEN_5526;
  assign _GEN_5528 = 9'h1cf == _T_82861 ? _T_70003 : _GEN_5527;
  assign _GEN_5529 = 9'h1d0 == _T_82861 ? _T_79643 : _GEN_5528;
  assign _GEN_5530 = 9'h1d1 == _T_82861 ? _T_71443 : _GEN_5529;
  assign _GEN_5531 = 9'h1d2 == _T_82861 ? _T_59843 : _GEN_5530;
  assign _GEN_5532 = 9'h1d3 == _T_82861 ? _T_49843 : _GEN_5531;
  assign _GEN_5533 = 9'h1d4 == _T_82861 ? _T_36003 : _GEN_5532;
  assign _GEN_5534 = 9'h1d5 == _T_82861 ? _T_81563 : _GEN_5533;
  assign _GEN_5535 = 9'h1d6 == _T_82861 ? _T_70323 : _GEN_5534;
  assign _GEN_5536 = 9'h1d7 == _T_82861 ? _T_53083 : _GEN_5535;
  assign _GEN_5537 = 9'h1d8 == _T_82861 ? _T_38723 : _GEN_5536;
  assign _GEN_5538 = 9'h1d9 == _T_82861 ? _T_66283 : _GEN_5537;
  assign _GEN_5539 = 9'h1da == _T_82861 ? _T_78683 : _GEN_5538;
  assign _GEN_5540 = 9'h1db == _T_82861 ? _T_42563 : _GEN_5539;
  assign _GEN_5541 = 9'h1dc == _T_82861 ? _T_53723 : _GEN_5540;
  assign _GEN_5542 = 9'h1dd == _T_82861 ? _T_62403 : _GEN_5541;
  assign _GEN_5543 = 9'h1de == _T_82861 ? _T_74683 : _GEN_5542;
  assign _GEN_5544 = 9'h1df == _T_82861 ? _T_35363 : _GEN_5543;
  assign _GEN_5545 = 9'h1e0 == _T_82861 ? _T_44163 : _GEN_5544;
  assign _GEN_5546 = 9'h1e1 == _T_82861 ? _T_36163 : _GEN_5545;
  assign _GEN_5547 = 9'h1e2 == _T_82861 ? _T_71923 : _GEN_5546;
  assign _GEN_5548 = 9'h1e3 == _T_82861 ? _T_63683 : _GEN_5547;
  assign _GEN_5549 = 9'h1e4 == _T_82861 ? _T_50003 : _GEN_5548;
  assign _GEN_5550 = 9'h1e5 == _T_82861 ? _T_43523 : _GEN_5549;
  assign _GEN_5551 = 9'h1e6 == _T_82861 ? _T_81243 : _GEN_5550;
  assign _GEN_5552 = 9'h1e7 == _T_82861 ? _T_67243 : _GEN_5551;
  assign _GEN_5553 = 9'h1e8 == _T_82861 ? _T_53403 : _GEN_5552;
  assign _GEN_5554 = 9'h1e9 == _T_82861 ? _T_54043 : _GEN_5553;
  assign _GEN_5555 = 9'h1ea == _T_82861 ? _T_66443 : _GEN_5554;
  assign _GEN_5556 = 9'h1eb == _T_82861 ? _T_82203 : _GEN_5555;
  assign _GEN_5557 = 9'h1ec == _T_82861 ? _T_42723 : _GEN_5556;
  assign _GEN_5558 = 9'h1ed == _T_82861 ? _T_51003 : _GEN_5557;
  assign _GEN_5559 = 9'h1ee == _T_82861 ? _T_62723 : _GEN_5558;
  assign _GEN_5560 = 9'h1ef == _T_82861 ? _T_72243 : _GEN_5559;
  assign _GEN_5561 = 9'h1f0 == _T_82861 ? _T_82523 : _GEN_5560;
  assign _GEN_5562 = 9'h1f1 == _T_82861 ? _T_71283 : _GEN_5561;
  assign _GEN_5563 = 9'h1f2 == _T_82861 ? _T_59683 : _GEN_5562;
  assign _GEN_5564 = 9'h1f3 == _T_82861 ? _T_52763 : _GEN_5563;
  assign _GEN_5565 = 9'h1f4 == _T_82861 ? _T_38563 : _GEN_5564;
  assign _GEN_5566 = 9'h1f5 == _T_82861 ? _T_80763 : _GEN_5565;
  assign _GEN_5567 = 9'h1f6 == _T_82861 ? _T_69843 : _GEN_5566;
  assign _GEN_5568 = 9'h1f7 == _T_82861 ? _T_55003 : _GEN_5567;
  assign _GEN_5569 = 9'h1f8 == _T_82861 ? _T_40483 : _GEN_5568;
  assign _GEN_5570 = 9'h1f9 == _T_82861 ? _T_65803 : _GEN_5569;
  assign _GEN_5571 = 9'h1fa == _T_82861 ? _T_78043 : _GEN_5570;
  assign _GEN_5572 = 9'h1fb == _T_82861 ? _T_45763 : _GEN_5571;
  assign _GEN_5573 = 9'h1fc == _T_82861 ? _T_55643 : _GEN_5572;
  assign _GEN_5574 = 9'h1fd == _T_82861 ? _T_61603 : _GEN_5573;
  assign _GEN_5575 = 9'h1fe == _T_82861 ? _T_74483 : _GEN_5574;
  assign _GEN_5576 = 9'h1ff == _T_82861 ? _T_37763 : _GEN_5575;
  assign _T_103419 = _GEN_5065 ? _GEN_5576 : 32'h0;
  assign _T_103420 = _T_25901[11:2];
  assign _T_103421 = _T_25901[1:0];
  assign _GEN_5577 = _T_1403 ? 8'h0 : _GEN_2460;
  assign _GEN_5578 = _T_1403 ? 8'h0 : _GEN_2461;
  assign _GEN_5579 = _T_1403 ? 8'h0 : _GEN_2462;
  assign _GEN_5580 = _T_1403 ? 8'h0 : _GEN_2463;
  assign _GEN_5581 = _T_1403 ? 8'h0 : _GEN_2473;
  assign _GEN_5582 = _T_1403 ? 8'h0 : _GEN_2474;
  assign _GEN_5583 = _T_1403 ? 8'h0 : _GEN_2475;
  assign _GEN_5584 = _T_1403 ? 8'h0 : _GEN_2476;
  assign _GEN_5585 = _T_1403 ? 8'h0 : _GEN_2486;
  assign _GEN_5586 = _T_1403 ? 8'h0 : _GEN_2487;
  assign _GEN_5587 = _T_1403 ? 8'h0 : _GEN_2488;
  assign _GEN_5588 = _T_1403 ? 8'h0 : _GEN_2489;
  assign _GEN_5589 = _T_1403 ? 8'h0 : _GEN_2499;
  assign _GEN_5590 = _T_1403 ? 8'h0 : _GEN_2500;
  assign _GEN_5591 = _T_1403 ? 8'h0 : _GEN_2501;
  assign _GEN_5592 = _T_1403 ? 8'h0 : _GEN_2502;
  assign _GEN_5593 = _T_1403 ? 8'h0 : _GEN_2447;
  assign _GEN_5594 = _T_1403 ? 8'h0 : _GEN_2448;
  assign _GEN_5595 = _T_1403 ? 8'h0 : _GEN_2449;
  assign _GEN_5596 = _T_1403 ? 8'h0 : _GEN_2450;
  assign _GEN_5597 = _T_1403 ? 8'h0 : _GEN_2464;
  assign _GEN_5598 = _T_1403 ? 8'h0 : _GEN_2465;
  assign _GEN_5599 = _T_1403 ? 8'h0 : _GEN_2466;
  assign _GEN_5600 = _T_1403 ? 8'h0 : _GEN_2467;
  assign _GEN_5601 = _T_1403 ? 8'h0 : _GEN_2477;
  assign _GEN_5602 = _T_1403 ? 8'h0 : _GEN_2478;
  assign _GEN_5603 = _T_1403 ? 8'h0 : _GEN_2479;
  assign _GEN_5604 = _T_1403 ? 8'h0 : _GEN_2480;
  assign _GEN_5605 = _T_1403 ? 8'h0 : _GEN_2495;
  assign _GEN_5606 = _T_1403 ? 8'h0 : _GEN_2496;
  assign _GEN_5607 = _T_1403 ? 8'h0 : _GEN_2497;
  assign _GEN_5608 = _T_1403 ? 8'h0 : _GEN_2498;
  assign _GEN_5609 = _T_1403 ? 8'h0 : _GEN_2503;
  assign _GEN_5610 = _T_1403 ? 8'h0 : _GEN_2504;
  assign _GEN_5611 = _T_1403 ? 8'h0 : _GEN_2505;
  assign _GEN_5612 = _T_1403 ? 8'h0 : _GEN_2506;
  assign _GEN_5613 = _T_1403 ? 8'h0 : _GEN_2443;
  assign _GEN_5614 = _T_1403 ? 8'h0 : _GEN_2444;
  assign _GEN_5615 = _T_1403 ? 8'h0 : _GEN_2445;
  assign _GEN_5616 = _T_1403 ? 8'h0 : _GEN_2446;
  assign _GEN_5617 = _T_1403 ? 8'h0 : _GEN_2439;
  assign _GEN_5618 = _T_1403 ? 8'h0 : _GEN_2440;
  assign _GEN_5619 = _T_1403 ? 8'h0 : _GEN_2441;
  assign _GEN_5620 = _T_1403 ? 8'h0 : _GEN_2442;
  assign _GEN_5621 = _T_1403 ? 8'h0 : _GEN_2491;
  assign _GEN_5622 = _T_1403 ? 8'h0 : _GEN_2492;
  assign _GEN_5623 = _T_1403 ? 8'h0 : _GEN_2493;
  assign _GEN_5624 = _T_1403 ? 8'h0 : _GEN_2494;
  assign _GEN_5625 = _T_1403 ? 8'h0 : _GEN_2469;
  assign _GEN_5626 = _T_1403 ? 8'h0 : _GEN_2470;
  assign _GEN_5627 = _T_1403 ? 8'h0 : _GEN_2471;
  assign _GEN_5628 = _T_1403 ? 8'h0 : _GEN_2472;
  assign _GEN_5629 = _T_1403 ? 8'h0 : _GEN_2455;
  assign _GEN_5630 = _T_1403 ? 8'h0 : _GEN_2456;
  assign _GEN_5631 = _T_1403 ? 8'h0 : _GEN_2457;
  assign _GEN_5632 = _T_1403 ? 8'h0 : _GEN_2458;
  assign _GEN_5633 = _T_1403 ? 8'h0 : _GEN_2451;
  assign _GEN_5634 = _T_1403 ? 8'h0 : _GEN_2452;
  assign _GEN_5635 = _T_1403 ? 8'h0 : _GEN_2453;
  assign _GEN_5636 = _T_1403 ? 8'h0 : _GEN_2454;
  assign _GEN_5637 = _T_1403 ? 8'h0 : _GEN_2507;
  assign _GEN_5638 = _T_1403 ? 8'h0 : _GEN_2508;
  assign _GEN_5639 = _T_1403 ? 8'h0 : _GEN_2509;
  assign _GEN_5640 = _T_1403 ? 8'h0 : _GEN_2510;
  assign _GEN_5641 = _T_1403 ? 8'h0 : _GEN_2482;
  assign _GEN_5642 = _T_1403 ? 8'h0 : _GEN_2483;
  assign _GEN_5643 = _T_1403 ? 8'h0 : _GEN_2484;
  assign _GEN_5644 = _T_1403 ? 8'h0 : _GEN_2485;
  assign _T_103511 = ctrlStateReg != 2'h0;
  assign _T_103513 = ctrlStateReg == 2'h0;
  assign _T_103515 = ctrlStateReg == 2'h0;
  assign _T_103517 = ctrlStateReg == 2'h0;
  assign _T_103519 = ctrlStateReg == 2'h0;
  assign _T_103521 = ctrlStateReg == 2'h0;
  assign _T_103522 = ~ _T_103513;
  assign _T_103523 = _T_5158 & _T_103522;
  assign _T_103525 = _T_3758 & _T_103522;
  assign _T_103526 = _T_103523 | _T_103525;
  assign _T_103528 = _T_6038 & _T_103522;
  assign _T_103529 = _T_103526 | _T_103528;
  assign _T_103531 = dmiAbstractDataAccess & _T_103522;
  assign _T_103532 = _T_103529 | _T_103531;
  assign _T_103534 = dmiProgramBufferAccess & _T_103522;
  assign _T_103535 = _T_103532 | _T_103534;
  assign commandWrIsAccessRegister = _T_2335 == 8'h0;
  assign commandRegIsAccessRegister = COMMANDRdData_cmdtype == 8'h0;
  assign _T_103539 = commandWrIsAccessRegister == 1'h0;
  assign commandWrIsUnsupported = COMMANDWrEn & _T_103539;
  assign _T_103545 = _T_23656 == 1'h0;
  assign _T_103547 = _T_23654 >= 16'h1000;
  assign _T_103549 = _T_23654 <= 16'h101f;
  assign _T_103550 = _T_103547 & _T_103549;
  assign _T_103551 = _T_103545 | _T_103550;
  assign _T_103553 = ~ haltedBitRegs_0;
  assign _GEN_5645 = _T_103551 ? 1'h0 : 1'h1;
  assign _GEN_5646 = _T_103551 ? _T_103553 : 1'h0;
  assign _GEN_5647 = commandRegIsAccessRegister ? _GEN_5645 : 1'h1;
  assign _GEN_5648 = commandRegIsAccessRegister ? _GEN_5646 : 1'h0;
  assign _T_103554 = COMMANDWrEn & commandWrIsAccessRegister;
  assign _T_103556 = ABSTRACTCSReg_cmderr == 3'h0;
  assign wrAccessRegisterCommand = _T_103554 & _T_103556;
  assign _T_103557 = autoexec & commandRegIsAccessRegister;
  assign regAccessRegisterCommand = _T_103557 & _T_103556;
  assign _T_103562 = wrAccessRegisterCommand | regAccessRegisterCommand;
  assign _GEN_5649 = _T_103562 ? 2'h1 : ctrlStateReg;
  assign _T_103565 = _T_103562 == 1'h0;
  assign _T_103566 = _T_103565 & commandWrIsUnsupported;
  assign _T_103568 = autoexec & _GEN_5647;
  assign _T_103572 = commandWrIsUnsupported == 1'h0;
  assign _T_103573 = _T_103565 & _T_103572;
  assign _T_103574 = _T_103573 & _T_103568;
  assign _GEN_5651 = _T_103574 ? 1'h1 : _T_103566;
  assign _GEN_5652 = _T_103513 ? _GEN_5649 : ctrlStateReg;
  assign _GEN_5653 = _T_103513 ? _GEN_5651 : 1'h0;
  assign _T_103577 = ctrlStateReg == 2'h1;
  assign _T_103579 = _T_103513 == 1'h0;
  assign _T_103580 = _T_103579 & _T_103577;
  assign _GEN_5654 = _GEN_5647 ? 1'h1 : _GEN_5653;
  assign _GEN_5655 = _GEN_5647 ? 2'h0 : _GEN_5652;
  assign _T_103584 = _GEN_5647 == 1'h0;
  assign _T_103585 = _T_103584 & _GEN_5648;
  assign _GEN_5657 = _T_103585 ? 2'h0 : _GEN_5655;
  assign _T_103591 = _GEN_5648 == 1'h0;
  assign _T_103592 = _T_103584 & _T_103591;
  assign _GEN_5658 = _T_103592 ? 2'h2 : _GEN_5657;
  assign _GEN_5660 = _T_103580 ? _GEN_5654 : _GEN_5653;
  assign _GEN_5661 = _T_103580 ? _GEN_5658 : _GEN_5652;
  assign _GEN_5662 = _T_103580 ? _T_103585 : 1'h0;
  assign _GEN_5663 = _T_103580 ? _T_103592 : 1'h0;
  assign _T_103596 = ctrlStateReg == 2'h2;
  assign _T_103600 = _T_103577 == 1'h0;
  assign _T_103601 = _T_103579 & _T_103600;
  assign _T_103602 = _T_103601 & _T_103596;
  assign _T_103604 = goReg == 1'h0;
  assign _T_103605 = _T_103604 & _T_57263;
  assign _T_103606 = _T_50184 == selectedHartReg;
  assign _T_103607 = _T_103605 & _T_103606;
  assign _GEN_5664 = _T_103607 ? 2'h0 : _GEN_5661;
  assign _GEN_5665 = _T_69183 ? 2'h0 : _GEN_5664;
  assign _GEN_5667 = _T_103602 ? _GEN_5665 : _GEN_5661;
  assign _GEN_5668 = _T_103602 ? _T_69183 : 1'h0;
  assign _GEN_5669 = _T_1403 ? 2'h0 : ctrlStateReg;
  assign _GEN_5670 = _T_1405 ? _GEN_5667 : _GEN_5669;
  assign _GEN_7411 = _T_1405 & _T_8236;
  assign _GEN_7413 = _T_103602 & _T_69183;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  haltedBitRegs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  resumeReqRegs_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  selectedHartReg = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  ABSTRACTCSReg_reserved0 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  ABSTRACTCSReg_progsize = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  ABSTRACTCSReg_reserved1 = _RAND_5[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  ABSTRACTCSReg_reserved2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  ABSTRACTCSReg_cmderr = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  ABSTRACTCSReg_reserved3 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  ABSTRACTCSReg_datacount = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  ABSTRACTAUTOReg_autoexecprogbuf = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  ABSTRACTAUTOReg_reserved0 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  ABSTRACTAUTOReg_autoexecdata = _RAND_12[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  COMMANDRdData_cmdtype = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  COMMANDRdData_control = _RAND_14[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  abstractDataMem_0 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  abstractDataMem_1 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  abstractDataMem_2 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  abstractDataMem_3 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  programBufferMem_0 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  programBufferMem_1 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  programBufferMem_2 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  programBufferMem_3 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  programBufferMem_4 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  programBufferMem_5 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  programBufferMem_6 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  programBufferMem_7 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  programBufferMem_8 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  programBufferMem_9 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  programBufferMem_10 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  programBufferMem_11 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  programBufferMem_12 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  programBufferMem_13 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  programBufferMem_14 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  programBufferMem_15 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  programBufferMem_16 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  programBufferMem_17 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  programBufferMem_18 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  programBufferMem_19 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  programBufferMem_20 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  programBufferMem_21 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  programBufferMem_22 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  programBufferMem_23 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  programBufferMem_24 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  programBufferMem_25 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  programBufferMem_26 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  programBufferMem_27 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  programBufferMem_28 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  programBufferMem_29 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  programBufferMem_30 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  programBufferMem_31 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  programBufferMem_32 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  programBufferMem_33 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  programBufferMem_34 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  programBufferMem_35 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  programBufferMem_36 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  programBufferMem_37 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  programBufferMem_38 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  programBufferMem_39 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  programBufferMem_40 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  programBufferMem_41 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  programBufferMem_42 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  programBufferMem_43 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  programBufferMem_44 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  programBufferMem_45 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  programBufferMem_46 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  programBufferMem_47 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  programBufferMem_48 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  programBufferMem_49 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  programBufferMem_50 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  programBufferMem_51 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  programBufferMem_52 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  programBufferMem_53 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  programBufferMem_54 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  programBufferMem_55 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  programBufferMem_56 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  programBufferMem_57 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  programBufferMem_58 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  programBufferMem_59 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  programBufferMem_60 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  programBufferMem_61 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  programBufferMem_62 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  programBufferMem_63 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  goReg = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  abstractGeneratedMem_0 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  abstractGeneratedMem_1 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  ctrlStateReg = _RAND_86[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      haltedBitRegs_0 <= 1'h0;
    end else begin
      if (_T_1405) begin
        if (_T_2790) begin
          if (_T_2792) begin
            haltedBitRegs_0 <= 1'h0;
          end else begin
            if (_T_57263) begin
              if (_T_2786) begin
                haltedBitRegs_0 <= 1'h1;
              end else begin
                if (_T_1403) begin
                  haltedBitRegs_0 <= 1'h0;
                end
              end
            end else begin
              if (_T_1403) begin
                haltedBitRegs_0 <= 1'h0;
              end
            end
          end
        end else begin
          if (_T_57263) begin
            if (_T_2786) begin
              haltedBitRegs_0 <= 1'h1;
            end else begin
              if (_T_1403) begin
                haltedBitRegs_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_1403) begin
              haltedBitRegs_0 <= 1'h0;
            end
          end
        end
      end else begin
        haltedBitRegs_0 <= _GEN_49;
      end
    end
    if (reset) begin
      resumeReqRegs_0 <= 1'h0;
    end else begin
      if (_T_1405) begin
        if (resumereq) begin
          resumeReqRegs_0 <= 1'h1;
        end else begin
          if (_T_63863) begin
            if (_T_2792) begin
              resumeReqRegs_0 <= 1'h0;
            end else begin
              if (_T_1403) begin
                resumeReqRegs_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_1403) begin
              resumeReqRegs_0 <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_1403) begin
          resumeReqRegs_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      selectedHartReg <= 10'h0;
    end else begin
      if (_T_1197) begin
        selectedHartReg <= io_innerCtrl_bits_hartsel;
      end
    end
    if (_T_1403) begin
      ABSTRACTCSReg_reserved0 <= 3'h0;
    end
    if (_T_1403) begin
      ABSTRACTCSReg_progsize <= 5'h10;
    end
    if (_T_1403) begin
      ABSTRACTCSReg_reserved1 <= 11'h0;
    end
    if (_T_1403) begin
      ABSTRACTCSReg_reserved2 <= 1'h0;
    end
    if (_T_1405) begin
      if (_T_1438) begin
        if (ABSTRACTCSWrEn) begin
          ABSTRACTCSReg_cmderr <= _T_1440;
        end else begin
          if (_T_1426) begin
            ABSTRACTCSReg_cmderr <= 3'h4;
          end else begin
            if (_T_1416) begin
              ABSTRACTCSReg_cmderr <= 3'h2;
            end else begin
              if (_T_1409) begin
                ABSTRACTCSReg_cmderr <= 3'h3;
              end else begin
                if (_T_103535) begin
                  ABSTRACTCSReg_cmderr <= 3'h1;
                end else begin
                  if (_T_1403) begin
                    ABSTRACTCSReg_cmderr <= 3'h0;
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_1426) begin
          ABSTRACTCSReg_cmderr <= 3'h4;
        end else begin
          if (_T_1416) begin
            ABSTRACTCSReg_cmderr <= 3'h2;
          end else begin
            if (_T_1409) begin
              ABSTRACTCSReg_cmderr <= 3'h3;
            end else begin
              if (_T_103535) begin
                ABSTRACTCSReg_cmderr <= 3'h1;
              end else begin
                if (_T_1403) begin
                  ABSTRACTCSReg_cmderr <= 3'h0;
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_1403) begin
        ABSTRACTCSReg_cmderr <= 3'h0;
      end
    end
    if (_T_1403) begin
      ABSTRACTCSReg_reserved3 <= 3'h0;
    end
    if (_T_1403) begin
      ABSTRACTCSReg_datacount <= 5'h1;
    end
    if (_T_1473) begin
      ABSTRACTAUTOReg_autoexecprogbuf <= _T_1462;
    end else begin
      if (_T_1403) begin
        ABSTRACTAUTOReg_autoexecprogbuf <= 16'h0;
      end
    end
    if (_T_1403) begin
      ABSTRACTAUTOReg_reserved0 <= 4'h0;
    end
    if (_T_1473) begin
      ABSTRACTAUTOReg_autoexecdata <= _T_1477;
    end else begin
      if (_T_1403) begin
        ABSTRACTAUTOReg_autoexecdata <= 12'h0;
      end
    end
    if (_T_1405) begin
      if (COMMANDWrEn) begin
        COMMANDRdData_cmdtype <= _T_2335;
      end else begin
        if (_T_1403) begin
          COMMANDRdData_cmdtype <= 8'h0;
        end
      end
    end else begin
      if (_T_1403) begin
        COMMANDRdData_cmdtype <= 8'h0;
      end
    end
    if (_T_1405) begin
      if (COMMANDWrEn) begin
        COMMANDRdData_control <= _T_2334;
      end else begin
        if (_T_1403) begin
          COMMANDRdData_control <= 24'h0;
        end
      end
    end else begin
      if (_T_1403) begin
        COMMANDRdData_control <= 24'h0;
      end
    end
    if (_T_1403) begin
      abstractDataMem_0 <= 8'h0;
    end else begin
      if (_T_51503) begin
        abstractDataMem_0 <= _T_35064;
      end else begin
        if (_T_7956) begin
          if (_T_6278) begin
            abstractDataMem_0 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      abstractDataMem_1 <= 8'h0;
    end else begin
      if (_T_51543) begin
        abstractDataMem_1 <= _T_35104;
      end else begin
        if (_T_7957) begin
          if (_T_6318) begin
            abstractDataMem_1 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      abstractDataMem_2 <= 8'h0;
    end else begin
      if (_T_51583) begin
        abstractDataMem_2 <= _T_35144;
      end else begin
        if (_T_7958) begin
          if (_T_6358) begin
            abstractDataMem_2 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      abstractDataMem_3 <= 8'h0;
    end else begin
      if (_T_51623) begin
        abstractDataMem_3 <= _T_35184;
      end else begin
        if (_T_7959) begin
          if (_T_6398) begin
            abstractDataMem_3 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_0 <= 8'h0;
    end else begin
      if (_T_62103) begin
        programBufferMem_0 <= _T_35064;
      end else begin
        if (_T_7960) begin
          if (_T_4598) begin
            programBufferMem_0 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_1 <= 8'h0;
    end else begin
      if (_T_62143) begin
        programBufferMem_1 <= _T_35104;
      end else begin
        if (_T_7961) begin
          if (_T_4638) begin
            programBufferMem_1 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_2 <= 8'h0;
    end else begin
      if (_T_62183) begin
        programBufferMem_2 <= _T_35144;
      end else begin
        if (_T_7962) begin
          if (_T_4678) begin
            programBufferMem_2 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_3 <= 8'h0;
    end else begin
      if (_T_62223) begin
        programBufferMem_3 <= _T_35184;
      end else begin
        if (_T_7963) begin
          if (_T_4718) begin
            programBufferMem_3 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_4 <= 8'h0;
    end else begin
      if (_T_66943) begin
        programBufferMem_4 <= _T_35064;
      end else begin
        if (_T_7964) begin
          if (_T_4278) begin
            programBufferMem_4 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_5 <= 8'h0;
    end else begin
      if (_T_66983) begin
        programBufferMem_5 <= _T_35104;
      end else begin
        if (_T_7965) begin
          if (_T_4318) begin
            programBufferMem_5 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_6 <= 8'h0;
    end else begin
      if (_T_67023) begin
        programBufferMem_6 <= _T_35144;
      end else begin
        if (_T_7966) begin
          if (_T_4358) begin
            programBufferMem_6 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_7 <= 8'h0;
    end else begin
      if (_T_67063) begin
        programBufferMem_7 <= _T_35184;
      end else begin
        if (_T_7967) begin
          if (_T_4398) begin
            programBufferMem_7 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_8 <= 8'h0;
    end else begin
      if (_T_77263) begin
        programBufferMem_8 <= _T_35064;
      end else begin
        if (_T_7968) begin
          if (_T_4758) begin
            programBufferMem_8 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_9 <= 8'h0;
    end else begin
      if (_T_77303) begin
        programBufferMem_9 <= _T_35104;
      end else begin
        if (_T_7969) begin
          if (_T_4798) begin
            programBufferMem_9 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_10 <= 8'h0;
    end else begin
      if (_T_77343) begin
        programBufferMem_10 <= _T_35144;
      end else begin
        if (_T_7970) begin
          if (_T_4838) begin
            programBufferMem_10 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_11 <= 8'h0;
    end else begin
      if (_T_77383) begin
        programBufferMem_11 <= _T_35184;
      end else begin
        if (_T_7971) begin
          if (_T_4878) begin
            programBufferMem_11 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_12 <= 8'h0;
    end else begin
      if (_T_43223) begin
        programBufferMem_12 <= _T_35064;
      end else begin
        if (_T_7972) begin
          if (_T_5518) begin
            programBufferMem_12 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_13 <= 8'h0;
    end else begin
      if (_T_43263) begin
        programBufferMem_13 <= _T_35104;
      end else begin
        if (_T_7973) begin
          if (_T_5558) begin
            programBufferMem_13 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_14 <= 8'h0;
    end else begin
      if (_T_43303) begin
        programBufferMem_14 <= _T_35144;
      end else begin
        if (_T_7974) begin
          if (_T_5598) begin
            programBufferMem_14 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_15 <= 8'h0;
    end else begin
      if (_T_43343) begin
        programBufferMem_15 <= _T_35184;
      end else begin
        if (_T_7975) begin
          if (_T_5638) begin
            programBufferMem_15 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_16 <= 8'h0;
    end else begin
      if (_T_54063) begin
        programBufferMem_16 <= _T_35064;
      end else begin
        if (_T_7976) begin
          if (_T_6078) begin
            programBufferMem_16 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_17 <= 8'h0;
    end else begin
      if (_T_54103) begin
        programBufferMem_17 <= _T_35104;
      end else begin
        if (_T_7977) begin
          if (_T_6118) begin
            programBufferMem_17 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_18 <= 8'h0;
    end else begin
      if (_T_54143) begin
        programBufferMem_18 <= _T_35144;
      end else begin
        if (_T_7978) begin
          if (_T_6158) begin
            programBufferMem_18 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_19 <= 8'h0;
    end else begin
      if (_T_54183) begin
        programBufferMem_19 <= _T_35184;
      end else begin
        if (_T_7979) begin
          if (_T_6198) begin
            programBufferMem_19 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_20 <= 8'h0;
    end else begin
      if (_T_63383) begin
        programBufferMem_20 <= _T_35064;
      end else begin
        if (_T_7980) begin
          if (_T_3798) begin
            programBufferMem_20 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_21 <= 8'h0;
    end else begin
      if (_T_63423) begin
        programBufferMem_21 <= _T_35104;
      end else begin
        if (_T_7981) begin
          if (_T_3838) begin
            programBufferMem_21 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_22 <= 8'h0;
    end else begin
      if (_T_63463) begin
        programBufferMem_22 <= _T_35144;
      end else begin
        if (_T_7982) begin
          if (_T_3878) begin
            programBufferMem_22 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_23 <= 8'h0;
    end else begin
      if (_T_63503) begin
        programBufferMem_23 <= _T_35184;
      end else begin
        if (_T_7983) begin
          if (_T_3918) begin
            programBufferMem_23 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_24 <= 8'h0;
    end else begin
      if (_T_75183) begin
        programBufferMem_24 <= _T_35064;
      end else begin
        if (_T_7984) begin
          if (_T_4118) begin
            programBufferMem_24 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_25 <= 8'h0;
    end else begin
      if (_T_75223) begin
        programBufferMem_25 <= _T_35104;
      end else begin
        if (_T_7985) begin
          if (_T_4158) begin
            programBufferMem_25 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_26 <= 8'h0;
    end else begin
      if (_T_75263) begin
        programBufferMem_26 <= _T_35144;
      end else begin
        if (_T_7986) begin
          if (_T_4198) begin
            programBufferMem_26 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_27 <= 8'h0;
    end else begin
      if (_T_75303) begin
        programBufferMem_27 <= _T_35184;
      end else begin
        if (_T_7987) begin
          if (_T_4238) begin
            programBufferMem_27 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_28 <= 8'h0;
    end else begin
      if (_T_81903) begin
        programBufferMem_28 <= _T_35064;
      end else begin
        if (_T_7988) begin
          if (_T_5358) begin
            programBufferMem_28 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_29 <= 8'h0;
    end else begin
      if (_T_81943) begin
        programBufferMem_29 <= _T_35104;
      end else begin
        if (_T_7989) begin
          if (_T_5398) begin
            programBufferMem_29 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_30 <= 8'h0;
    end else begin
      if (_T_81983) begin
        programBufferMem_30 <= _T_35144;
      end else begin
        if (_T_7990) begin
          if (_T_5438) begin
            programBufferMem_30 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_31 <= 8'h0;
    end else begin
      if (_T_82023) begin
        programBufferMem_31 <= _T_35184;
      end else begin
        if (_T_7991) begin
          if (_T_5478) begin
            programBufferMem_31 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_32 <= 8'h0;
    end else begin
      if (_T_42263) begin
        programBufferMem_32 <= _T_35064;
      end else begin
        if (_T_7992) begin
          if (_T_5878) begin
            programBufferMem_32 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_33 <= 8'h0;
    end else begin
      if (_T_42303) begin
        programBufferMem_33 <= _T_35104;
      end else begin
        if (_T_7993) begin
          if (_T_5918) begin
            programBufferMem_33 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_34 <= 8'h0;
    end else begin
      if (_T_42343) begin
        programBufferMem_34 <= _T_35144;
      end else begin
        if (_T_7994) begin
          if (_T_5958) begin
            programBufferMem_34 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_35 <= 8'h0;
    end else begin
      if (_T_42383) begin
        programBufferMem_35 <= _T_35184;
      end else begin
        if (_T_7995) begin
          if (_T_5998) begin
            programBufferMem_35 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_36 <= 8'h0;
    end else begin
      if (_T_36663) begin
        programBufferMem_36 <= _T_35064;
      end else begin
        if (_T_7996) begin
          if (_T_4438) begin
            programBufferMem_36 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_37 <= 8'h0;
    end else begin
      if (_T_36703) begin
        programBufferMem_37 <= _T_35104;
      end else begin
        if (_T_7997) begin
          if (_T_4478) begin
            programBufferMem_37 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_38 <= 8'h0;
    end else begin
      if (_T_36743) begin
        programBufferMem_38 <= _T_35144;
      end else begin
        if (_T_7998) begin
          if (_T_4518) begin
            programBufferMem_38 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_39 <= 8'h0;
    end else begin
      if (_T_36783) begin
        programBufferMem_39 <= _T_35184;
      end else begin
        if (_T_7999) begin
          if (_T_4558) begin
            programBufferMem_39 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_40 <= 8'h0;
    end else begin
      if (_T_72263) begin
        programBufferMem_40 <= _T_35064;
      end else begin
        if (_T_8000) begin
          if (_T_3598) begin
            programBufferMem_40 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_41 <= 8'h0;
    end else begin
      if (_T_72303) begin
        programBufferMem_41 <= _T_35104;
      end else begin
        if (_T_8001) begin
          if (_T_3638) begin
            programBufferMem_41 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_42 <= 8'h0;
    end else begin
      if (_T_72343) begin
        programBufferMem_42 <= _T_35144;
      end else begin
        if (_T_8002) begin
          if (_T_3678) begin
            programBufferMem_42 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_43 <= 8'h0;
    end else begin
      if (_T_72383) begin
        programBufferMem_43 <= _T_35184;
      end else begin
        if (_T_8003) begin
          if (_T_3718) begin
            programBufferMem_43 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_44 <= 8'h0;
    end else begin
      if (_T_60343) begin
        programBufferMem_44 <= _T_35064;
      end else begin
        if (_T_8004) begin
          if (_T_5718) begin
            programBufferMem_44 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_45 <= 8'h0;
    end else begin
      if (_T_60383) begin
        programBufferMem_45 <= _T_35104;
      end else begin
        if (_T_8005) begin
          if (_T_5758) begin
            programBufferMem_45 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_46 <= 8'h0;
    end else begin
      if (_T_60423) begin
        programBufferMem_46 <= _T_35144;
      end else begin
        if (_T_8006) begin
          if (_T_5798) begin
            programBufferMem_46 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_47 <= 8'h0;
    end else begin
      if (_T_60463) begin
        programBufferMem_47 <= _T_35184;
      end else begin
        if (_T_8007) begin
          if (_T_5838) begin
            programBufferMem_47 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_48 <= 8'h0;
    end else begin
      if (_T_47583) begin
        programBufferMem_48 <= _T_35064;
      end else begin
        if (_T_8008) begin
          if (_T_5198) begin
            programBufferMem_48 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_49 <= 8'h0;
    end else begin
      if (_T_47623) begin
        programBufferMem_49 <= _T_35104;
      end else begin
        if (_T_8009) begin
          if (_T_5238) begin
            programBufferMem_49 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_50 <= 8'h0;
    end else begin
      if (_T_47663) begin
        programBufferMem_50 <= _T_35144;
      end else begin
        if (_T_8010) begin
          if (_T_5278) begin
            programBufferMem_50 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_51 <= 8'h0;
    end else begin
      if (_T_47703) begin
        programBufferMem_51 <= _T_35184;
      end else begin
        if (_T_8011) begin
          if (_T_5318) begin
            programBufferMem_51 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_52 <= 8'h0;
    end else begin
      if (_T_44503) begin
        programBufferMem_52 <= _T_35064;
      end else begin
        if (_T_8012) begin
          if (_T_4918) begin
            programBufferMem_52 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_53 <= 8'h0;
    end else begin
      if (_T_44543) begin
        programBufferMem_53 <= _T_35104;
      end else begin
        if (_T_8013) begin
          if (_T_4958) begin
            programBufferMem_53 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_54 <= 8'h0;
    end else begin
      if (_T_44583) begin
        programBufferMem_54 <= _T_35144;
      end else begin
        if (_T_8014) begin
          if (_T_4998) begin
            programBufferMem_54 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_55 <= 8'h0;
    end else begin
      if (_T_44623) begin
        programBufferMem_55 <= _T_35184;
      end else begin
        if (_T_8015) begin
          if (_T_5038) begin
            programBufferMem_55 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_56 <= 8'h0;
    end else begin
      if (_T_82223) begin
        programBufferMem_56 <= _T_35064;
      end else begin
        if (_T_8016) begin
          if (_T_3958) begin
            programBufferMem_56 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_57 <= 8'h0;
    end else begin
      if (_T_82263) begin
        programBufferMem_57 <= _T_35104;
      end else begin
        if (_T_8017) begin
          if (_T_3998) begin
            programBufferMem_57 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_58 <= 8'h0;
    end else begin
      if (_T_82303) begin
        programBufferMem_58 <= _T_35144;
      end else begin
        if (_T_8018) begin
          if (_T_4038) begin
            programBufferMem_58 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_59 <= 8'h0;
    end else begin
      if (_T_82343) begin
        programBufferMem_59 <= _T_35184;
      end else begin
        if (_T_8019) begin
          if (_T_4078) begin
            programBufferMem_59 <= _T_3719;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_60 <= 8'h0;
    end else begin
      if (_T_64863) begin
        programBufferMem_60 <= _T_35064;
      end else begin
        if (_T_8020) begin
          if (_T_6438) begin
            programBufferMem_60 <= _T_3599;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_61 <= 8'h0;
    end else begin
      if (_T_64903) begin
        programBufferMem_61 <= _T_35104;
      end else begin
        if (_T_8021) begin
          if (_T_6478) begin
            programBufferMem_61 <= _T_3639;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_62 <= 8'h0;
    end else begin
      if (_T_64943) begin
        programBufferMem_62 <= _T_35144;
      end else begin
        if (_T_8022) begin
          if (_T_6518) begin
            programBufferMem_62 <= _T_3679;
          end
        end
      end
    end
    if (_T_1403) begin
      programBufferMem_63 <= 8'h0;
    end else begin
      if (_T_64983) begin
        programBufferMem_63 <= _T_35184;
      end else begin
        if (_T_8023) begin
          if (_T_6558) begin
            programBufferMem_63 <= _T_3719;
          end
        end
      end
    end
    if (_T_1405) begin
      if (_T_8236) begin
        goReg <= 1'h0;
      end else begin
        if (_GEN_5663) begin
          goReg <= 1'h1;
        end else begin
          if (_T_1403) begin
            goReg <= 1'h0;
          end
        end
      end
    end else begin
      if (_T_1403) begin
        goReg <= 1'h0;
      end
    end
    if (_GEN_5663) begin
      if (_T_23656) begin
        if (_T_23655) begin
          abstractGeneratedMem_0 <= _T_23722;
        end else begin
          abstractGeneratedMem_0 <= _T_23727;
        end
      end else begin
        abstractGeneratedMem_0 <= 32'h13;
      end
    end
    if (_GEN_5663) begin
      if (_T_23657) begin
        abstractGeneratedMem_1 <= 32'h13;
      end else begin
        abstractGeneratedMem_1 <= 32'h100073;
      end
    end
    if (_T_1405) begin
      if (_T_103602) begin
        if (_T_69183) begin
          ctrlStateReg <= 2'h0;
        end else begin
          if (_T_103607) begin
            ctrlStateReg <= 2'h0;
          end else begin
            if (_T_103580) begin
              if (_T_103592) begin
                ctrlStateReg <= 2'h2;
              end else begin
                if (_T_103585) begin
                  ctrlStateReg <= 2'h0;
                end else begin
                  if (_GEN_5647) begin
                    ctrlStateReg <= 2'h0;
                  end else begin
                    if (_T_103513) begin
                      if (_T_103562) begin
                        ctrlStateReg <= 2'h1;
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_103513) begin
                if (_T_103562) begin
                  ctrlStateReg <= 2'h1;
                end
              end
            end
          end
        end
      end else begin
        if (_T_103580) begin
          if (_T_103592) begin
            ctrlStateReg <= 2'h2;
          end else begin
            if (_T_103585) begin
              ctrlStateReg <= 2'h0;
            end else begin
              if (_GEN_5647) begin
                ctrlStateReg <= 2'h0;
              end else begin
                if (_T_103513) begin
                  if (_T_103562) begin
                    ctrlStateReg <= 2'h1;
                  end
                end
              end
            end
          end
        end else begin
          if (_T_103513) begin
            if (_T_103562) begin
              ctrlStateReg <= 2'h1;
            end
          end
        end
      end
    end else begin
      if (_T_1403) begin
        ctrlStateReg <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7411 & _T_8241) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected 'GOING' hart.\n    at Debug.scala:767 assert(hartGoingId === 0.U, \"Unexpected 'GOING' hart.\")//Chisel3 #540 %%x, expected %%x\", hartGoingId, 0.U)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7411 & _T_8241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: HartSel to HartId Mapping is illegal for this Debug Implementation, because HartID must be < 1024 for it to work.\n    at Debug.scala:779 assert ((cfg.hartSelToHartId(selectedHartReg) < 1024.U),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7413 & _T_8241) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected 'EXCEPTION' hart\n    at Debug.scala:993 assert(hartExceptionId === 0.U, \"Unexpected 'EXCEPTION' hart\")//Chisel3 #540, %%x, expected %%x\", hartExceptionId, 0.U)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7413 & _T_8241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AsyncQueueSink_1(
  input         clock,
  input         reset,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_size,
  output        io_deq_bits_source,
  output [8:0]  io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data,
  output        io_ridx,
  input         io_widx,
  input  [2:0]  io_mem_0_opcode,
  input  [1:0]  io_mem_0_size,
  input         io_mem_0_source,
  input  [8:0]  io_mem_0_address,
  input  [3:0]  io_mem_0_mask,
  input  [31:0] io_mem_0_data,
  input         io_source_reset_n,
  output        io_ridx_valid,
  input         io_widx_valid
);
  wire  source_ready;
  wire  _T_17;
  wire  _T_19;
  wire  ridx_bin_clock;
  wire  ridx_bin_reset;
  wire  ridx_bin_io_d;
  wire  ridx_bin_io_q;
  wire  ridx_bin_io_en;
  wire [1:0] _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_28;
  wire  ridx;
  wire  widx_gray_sync_0_clock;
  wire  widx_gray_sync_0_reset;
  wire  widx_gray_sync_0_io_d;
  wire  widx_gray_sync_0_io_q;
  wire  widx_gray_sync_0_io_en;
  wire  widx_gray_sync_1_clock;
  wire  widx_gray_sync_1_reset;
  wire  widx_gray_sync_1_io_d;
  wire  widx_gray_sync_1_io_q;
  wire  widx_gray_sync_1_io_en;
  wire  widx_gray_sync_2_clock;
  wire  widx_gray_sync_2_reset;
  wire  widx_gray_sync_2_io_d;
  wire  widx_gray_sync_2_io_q;
  wire  widx_gray_sync_2_io_en;
  wire  _T_32;
  wire  valid;
  reg [2:0] _T_36_opcode;
  reg [31:0] _RAND_0;
  reg [1:0] _T_36_size;
  reg [31:0] _RAND_1;
  reg  _T_36_source;
  reg [31:0] _RAND_2;
  reg [8:0] _T_36_address;
  reg [31:0] _RAND_3;
  reg [3:0] _T_36_mask;
  reg [31:0] _RAND_4;
  reg [31:0] _T_36_data;
  reg [31:0] _RAND_5;
  wire [2:0] _GEN_0;
  wire [1:0] _GEN_2;
  wire  _GEN_3;
  wire [8:0] _GEN_4;
  wire [3:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire  valid_reg_clock;
  wire  valid_reg_reset;
  wire  valid_reg_io_d;
  wire  valid_reg_io_q;
  wire  valid_reg_io_en;
  wire  valid_reg_1;
  wire  _T_38;
  wire  ridx_gray_clock;
  wire  ridx_gray_reset;
  wire  ridx_gray_io_d;
  wire  ridx_gray_io_q;
  wire  ridx_gray_io_en;
  wire  AsyncValidSync_clock;
  wire  AsyncValidSync_reset;
  wire  AsyncValidSync_io_in;
  wire  AsyncValidSync_io_out;
  wire  AsyncValidSync_1_clock;
  wire  AsyncValidSync_1_reset;
  wire  AsyncValidSync_1_io_in;
  wire  AsyncValidSync_1_io_out;
  wire  AsyncValidSync_2_clock;
  wire  AsyncValidSync_2_reset;
  wire  AsyncValidSync_2_io_in;
  wire  AsyncValidSync_2_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  _T_60;
  wire  AsyncResetRegVec_clock;
  wire  AsyncResetRegVec_reset;
  wire  AsyncResetRegVec_io_d;
  wire  AsyncResetRegVec_io_q;
  wire  AsyncResetRegVec_io_en;
  AsyncResetRegVec_1 ridx_bin (
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_0 (
    .clock(widx_gray_sync_0_clock),
    .reset(widx_gray_sync_0_reset),
    .io_d(widx_gray_sync_0_io_d),
    .io_q(widx_gray_sync_0_io_q),
    .io_en(widx_gray_sync_0_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_1 (
    .clock(widx_gray_sync_1_clock),
    .reset(widx_gray_sync_1_reset),
    .io_d(widx_gray_sync_1_io_d),
    .io_q(widx_gray_sync_1_io_q),
    .io_en(widx_gray_sync_1_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_2 (
    .clock(widx_gray_sync_2_clock),
    .reset(widx_gray_sync_2_reset),
    .io_d(widx_gray_sync_2_io_d),
    .io_q(widx_gray_sync_2_io_q),
    .io_en(widx_gray_sync_2_io_en)
  );
  AsyncResetRegVec_1 valid_reg (
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_1 ridx_gray (
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync_3 AsyncValidSync (
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_4 AsyncValidSync_1 (
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_5 AsyncValidSync_2 (
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_1 AsyncResetRegVec (
    .clock(AsyncResetRegVec_clock),
    .reset(AsyncResetRegVec_reset),
    .io_d(AsyncResetRegVec_io_d),
    .io_q(AsyncResetRegVec_io_q),
    .io_en(AsyncResetRegVec_io_en)
  );
  assign io_deq_valid = _T_38;
  assign io_deq_bits_opcode = _T_36_opcode;
  assign io_deq_bits_size = _T_36_size;
  assign io_deq_bits_source = _T_36_source;
  assign io_deq_bits_address = _T_36_address;
  assign io_deq_bits_mask = _T_36_mask;
  assign io_deq_bits_data = _T_36_data;
  assign io_ridx = ridx_gray_io_q;
  assign io_ridx_valid = AsyncValidSync_io_out;
  assign source_ready = AsyncValidSync_2_io_out;
  assign _T_17 = io_deq_ready & io_deq_valid;
  assign _T_19 = source_ready == 1'h0;
  assign ridx_bin_clock = clock;
  assign ridx_bin_reset = reset;
  assign ridx_bin_io_d = _T_26;
  assign ridx_bin_io_en = 1'h1;
  assign _T_24 = ridx_bin_io_q + _T_17;
  assign _T_25 = _T_24[0:0];
  assign _T_26 = _T_19 ? 1'h0 : _T_25;
  assign _T_28 = _T_26 >> 1'h1;
  assign ridx = _T_26 ^ _T_28;
  assign widx_gray_sync_0_clock = clock;
  assign widx_gray_sync_0_reset = reset;
  assign widx_gray_sync_0_io_d = widx_gray_sync_1_io_q;
  assign widx_gray_sync_0_io_en = 1'h1;
  assign widx_gray_sync_1_clock = clock;
  assign widx_gray_sync_1_reset = reset;
  assign widx_gray_sync_1_io_d = widx_gray_sync_2_io_q;
  assign widx_gray_sync_1_io_en = 1'h1;
  assign widx_gray_sync_2_clock = clock;
  assign widx_gray_sync_2_reset = reset;
  assign widx_gray_sync_2_io_d = io_widx;
  assign widx_gray_sync_2_io_en = 1'h1;
  assign _T_32 = ridx != widx_gray_sync_0_io_q;
  assign valid = source_ready & _T_32;
  assign _GEN_0 = valid ? io_mem_0_opcode : _T_36_opcode;
  assign _GEN_2 = valid ? io_mem_0_size : _T_36_size;
  assign _GEN_3 = valid ? io_mem_0_source : _T_36_source;
  assign _GEN_4 = valid ? io_mem_0_address : _T_36_address;
  assign _GEN_5 = valid ? io_mem_0_mask : _T_36_mask;
  assign _GEN_6 = valid ? io_mem_0_data : _T_36_data;
  assign valid_reg_clock = clock;
  assign valid_reg_reset = reset;
  assign valid_reg_io_d = valid;
  assign valid_reg_io_en = 1'h1;
  assign valid_reg_1 = valid_reg_io_q;
  assign _T_38 = valid_reg_1 & source_ready;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = ridx;
  assign ridx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_43;
  assign AsyncValidSync_io_in = 1'h1;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_43;
  assign AsyncValidSync_1_io_in = io_widx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign _T_42 = io_source_reset_n == 1'h0;
  assign _T_43 = reset | _T_42;
  assign _T_60 = io_widx == io_ridx;
  assign AsyncResetRegVec_clock = clock;
  assign AsyncResetRegVec_reset = reset;
  assign AsyncResetRegVec_io_d = _T_60;
  assign AsyncResetRegVec_io_en = 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_36_opcode = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_36_size = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_36_source = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_36_address = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_36_mask = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_36_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (valid) begin
      _T_36_opcode <= io_mem_0_opcode;
    end
    if (valid) begin
      _T_36_size <= io_mem_0_size;
    end
    if (valid) begin
      _T_36_source <= io_mem_0_source;
    end
    if (valid) begin
      _T_36_address <= io_mem_0_address;
    end
    if (valid) begin
      _T_36_mask <= io_mem_0_mask;
    end
    if (valid) begin
      _T_36_data <= io_mem_0_data;
    end
  end
endmodule
module AsyncQueueSource_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [1:0]  io_enq_bits_size,
  input         io_enq_bits_source,
  input         io_enq_bits_sink,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_ridx,
  output        io_widx,
  output [2:0]  io_mem_0_opcode,
  output [1:0]  io_mem_0_param,
  output [1:0]  io_mem_0_size,
  output        io_mem_0_source,
  output        io_mem_0_sink,
  output [31:0] io_mem_0_data,
  output        io_mem_0_error,
  input         io_sink_reset_n,
  input         io_ridx_valid,
  output        io_widx_valid
);
  wire  sink_ready;
  reg [2:0] mem_0_opcode;
  reg [31:0] _RAND_0;
  reg [1:0] mem_0_param;
  reg [31:0] _RAND_1;
  reg [1:0] mem_0_size;
  reg [31:0] _RAND_2;
  reg  mem_0_source;
  reg [31:0] _RAND_3;
  reg  mem_0_sink;
  reg [31:0] _RAND_4;
  reg [31:0] mem_0_data;
  reg [31:0] _RAND_5;
  reg  mem_0_error;
  reg [31:0] _RAND_6;
  wire  _T_26;
  wire  _T_28;
  wire  widx_bin_clock;
  wire  widx_bin_reset;
  wire  widx_bin_io_d;
  wire  widx_bin_io_q;
  wire  widx_bin_io_en;
  wire [1:0] _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_37;
  wire  widx;
  wire  ridx_gray_sync_0_clock;
  wire  ridx_gray_sync_0_reset;
  wire  ridx_gray_sync_0_io_d;
  wire  ridx_gray_sync_0_io_q;
  wire  ridx_gray_sync_0_io_en;
  wire  ridx_gray_sync_1_clock;
  wire  ridx_gray_sync_1_reset;
  wire  ridx_gray_sync_1_io_d;
  wire  ridx_gray_sync_1_io_q;
  wire  ridx_gray_sync_1_io_en;
  wire  ridx_gray_sync_2_clock;
  wire  ridx_gray_sync_2_reset;
  wire  ridx_gray_sync_2_io_d;
  wire  ridx_gray_sync_2_io_q;
  wire  ridx_gray_sync_2_io_en;
  wire  _T_42;
  wire  _T_43;
  wire  ready;
  wire [2:0] _GEN_0;
  wire [1:0] _GEN_1;
  wire [1:0] _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [31:0] _GEN_5;
  wire  _GEN_6;
  wire  ready_reg_clock;
  wire  ready_reg_reset;
  wire  ready_reg_io_d;
  wire  ready_reg_io_q;
  wire  ready_reg_io_en;
  wire  ready_reg_1;
  wire  _T_48;
  wire  widx_gray_clock;
  wire  widx_gray_reset;
  wire  widx_gray_io_d;
  wire  widx_gray_io_q;
  wire  widx_gray_io_en;
  wire  AsyncValidSync_clock;
  wire  AsyncValidSync_reset;
  wire  AsyncValidSync_io_in;
  wire  AsyncValidSync_io_out;
  wire  AsyncValidSync_1_clock;
  wire  AsyncValidSync_1_reset;
  wire  AsyncValidSync_1_io_in;
  wire  AsyncValidSync_1_io_out;
  wire  AsyncValidSync_2_clock;
  wire  AsyncValidSync_2_reset;
  wire  AsyncValidSync_2_io_in;
  wire  AsyncValidSync_2_io_out;
  wire  _T_52;
  wire  _T_53;
  AsyncResetRegVec_1 widx_bin (
    .clock(widx_bin_clock),
    .reset(widx_bin_reset),
    .io_d(widx_bin_io_d),
    .io_q(widx_bin_io_q),
    .io_en(widx_bin_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_0 (
    .clock(ridx_gray_sync_0_clock),
    .reset(ridx_gray_sync_0_reset),
    .io_d(ridx_gray_sync_0_io_d),
    .io_q(ridx_gray_sync_0_io_q),
    .io_en(ridx_gray_sync_0_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_1 (
    .clock(ridx_gray_sync_1_clock),
    .reset(ridx_gray_sync_1_reset),
    .io_d(ridx_gray_sync_1_io_d),
    .io_q(ridx_gray_sync_1_io_q),
    .io_en(ridx_gray_sync_1_io_en)
  );
  AsyncResetRegVec_1 ridx_gray_sync_2 (
    .clock(ridx_gray_sync_2_clock),
    .reset(ridx_gray_sync_2_reset),
    .io_d(ridx_gray_sync_2_io_d),
    .io_q(ridx_gray_sync_2_io_q),
    .io_en(ridx_gray_sync_2_io_en)
  );
  AsyncResetRegVec_1 ready_reg (
    .clock(ready_reg_clock),
    .reset(ready_reg_reset),
    .io_d(ready_reg_io_d),
    .io_q(ready_reg_io_q),
    .io_en(ready_reg_io_en)
  );
  AsyncResetRegVec_1 widx_gray (
    .clock(widx_gray_clock),
    .reset(widx_gray_reset),
    .io_d(widx_gray_io_d),
    .io_q(widx_gray_io_q),
    .io_en(widx_gray_io_en)
  );
  AsyncValidSync AsyncValidSync (
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_1 AsyncValidSync_1 (
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_2 AsyncValidSync_2 (
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  assign io_enq_ready = _T_48;
  assign io_widx = widx_gray_io_q;
  assign io_mem_0_opcode = mem_0_opcode;
  assign io_mem_0_param = mem_0_param;
  assign io_mem_0_size = mem_0_size;
  assign io_mem_0_source = mem_0_source;
  assign io_mem_0_sink = mem_0_sink;
  assign io_mem_0_data = mem_0_data;
  assign io_mem_0_error = mem_0_error;
  assign io_widx_valid = AsyncValidSync_io_out;
  assign sink_ready = AsyncValidSync_2_io_out;
  assign _T_26 = io_enq_ready & io_enq_valid;
  assign _T_28 = sink_ready == 1'h0;
  assign widx_bin_clock = clock;
  assign widx_bin_reset = reset;
  assign widx_bin_io_d = _T_35;
  assign widx_bin_io_en = 1'h1;
  assign _T_33 = widx_bin_io_q + _T_26;
  assign _T_34 = _T_33[0:0];
  assign _T_35 = _T_28 ? 1'h0 : _T_34;
  assign _T_37 = _T_35 >> 1'h1;
  assign widx = _T_35 ^ _T_37;
  assign ridx_gray_sync_0_clock = clock;
  assign ridx_gray_sync_0_reset = reset;
  assign ridx_gray_sync_0_io_d = ridx_gray_sync_1_io_q;
  assign ridx_gray_sync_0_io_en = 1'h1;
  assign ridx_gray_sync_1_clock = clock;
  assign ridx_gray_sync_1_reset = reset;
  assign ridx_gray_sync_1_io_d = ridx_gray_sync_2_io_q;
  assign ridx_gray_sync_1_io_en = 1'h1;
  assign ridx_gray_sync_2_clock = clock;
  assign ridx_gray_sync_2_reset = reset;
  assign ridx_gray_sync_2_io_d = io_ridx;
  assign ridx_gray_sync_2_io_en = 1'h1;
  assign _T_42 = ridx_gray_sync_0_io_q ^ 1'h1;
  assign _T_43 = widx != _T_42;
  assign ready = sink_ready & _T_43;
  assign _GEN_0 = _T_26 ? io_enq_bits_opcode : mem_0_opcode;
  assign _GEN_1 = _T_26 ? io_enq_bits_param : mem_0_param;
  assign _GEN_2 = _T_26 ? io_enq_bits_size : mem_0_size;
  assign _GEN_3 = _T_26 ? io_enq_bits_source : mem_0_source;
  assign _GEN_4 = _T_26 ? io_enq_bits_sink : mem_0_sink;
  assign _GEN_5 = _T_26 ? io_enq_bits_data : mem_0_data;
  assign _GEN_6 = _T_26 ? io_enq_bits_error : mem_0_error;
  assign ready_reg_clock = clock;
  assign ready_reg_reset = reset;
  assign ready_reg_io_d = ready;
  assign ready_reg_io_en = 1'h1;
  assign ready_reg_1 = ready_reg_io_q;
  assign _T_48 = ready_reg_1 & sink_ready;
  assign widx_gray_clock = clock;
  assign widx_gray_reset = reset;
  assign widx_gray_io_d = widx;
  assign widx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_53;
  assign AsyncValidSync_io_in = 1'h1;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_53;
  assign AsyncValidSync_1_io_in = io_ridx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign _T_52 = io_sink_reset_n == 1'h0;
  assign _T_53 = reset | _T_52;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  mem_0_opcode = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0_param = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem_0_size = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_0_source = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  mem_0_sink = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_0_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  mem_0_error = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_26) begin
      mem_0_opcode <= io_enq_bits_opcode;
    end
    if (_T_26) begin
      mem_0_param <= io_enq_bits_param;
    end
    if (_T_26) begin
      mem_0_size <= io_enq_bits_size;
    end
    if (_T_26) begin
      mem_0_source <= io_enq_bits_source;
    end
    if (_T_26) begin
      mem_0_sink <= io_enq_bits_sink;
    end
    if (_T_26) begin
      mem_0_data <= io_enq_bits_data;
    end
    if (_T_26) begin
      mem_0_error <= io_enq_bits_error;
    end
  end
endmodule
module TLAsyncCrossingSink(
  input         clock,
  input         reset,
  input  [2:0]  io_in_0_a_mem_0_opcode,
  input  [1:0]  io_in_0_a_mem_0_size,
  input         io_in_0_a_mem_0_source,
  input  [8:0]  io_in_0_a_mem_0_address,
  input  [3:0]  io_in_0_a_mem_0_mask,
  input  [31:0] io_in_0_a_mem_0_data,
  output        io_in_0_a_ridx,
  input         io_in_0_a_widx,
  output        io_in_0_a_ridx_valid,
  input         io_in_0_a_widx_valid,
  input         io_in_0_a_source_reset_n,
  output        io_in_0_a_sink_reset_n,
  output [2:0]  io_in_0_d_mem_0_opcode,
  output [1:0]  io_in_0_d_mem_0_param,
  output [1:0]  io_in_0_d_mem_0_size,
  output        io_in_0_d_mem_0_source,
  output        io_in_0_d_mem_0_sink,
  output [31:0] io_in_0_d_mem_0_data,
  output        io_in_0_d_mem_0_error,
  input         io_in_0_d_ridx,
  output        io_in_0_d_widx,
  input         io_in_0_d_ridx_valid,
  output        io_in_0_d_widx_valid,
  output        io_in_0_d_source_reset_n,
  input         io_in_0_d_sink_reset_n,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [1:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [8:0]  io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [1:0]  io_out_0_d_bits_size,
  input         io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  AsyncQueueSink_clock;
  wire  AsyncQueueSink_reset;
  wire  AsyncQueueSink_io_deq_ready;
  wire  AsyncQueueSink_io_deq_valid;
  wire [2:0] AsyncQueueSink_io_deq_bits_opcode;
  wire [1:0] AsyncQueueSink_io_deq_bits_size;
  wire  AsyncQueueSink_io_deq_bits_source;
  wire [8:0] AsyncQueueSink_io_deq_bits_address;
  wire [3:0] AsyncQueueSink_io_deq_bits_mask;
  wire [31:0] AsyncQueueSink_io_deq_bits_data;
  wire  AsyncQueueSink_io_ridx;
  wire  AsyncQueueSink_io_widx;
  wire [2:0] AsyncQueueSink_io_mem_0_opcode;
  wire [1:0] AsyncQueueSink_io_mem_0_size;
  wire  AsyncQueueSink_io_mem_0_source;
  wire [8:0] AsyncQueueSink_io_mem_0_address;
  wire [3:0] AsyncQueueSink_io_mem_0_mask;
  wire [31:0] AsyncQueueSink_io_mem_0_data;
  wire  AsyncQueueSink_io_source_reset_n;
  wire  AsyncQueueSink_io_ridx_valid;
  wire  AsyncQueueSink_io_widx_valid;
  wire  _T_105;
  wire  _T_110_valid;
  wire [2:0] _T_110_bits_opcode;
  wire [1:0] _T_110_bits_size;
  wire  _T_110_bits_source;
  wire [8:0] _T_110_bits_address;
  wire [3:0] _T_110_bits_mask;
  wire [31:0] _T_110_bits_data;
  wire  AsyncQueueSource_clock;
  wire  AsyncQueueSource_reset;
  wire  AsyncQueueSource_io_enq_ready;
  wire  AsyncQueueSource_io_enq_valid;
  wire [2:0] AsyncQueueSource_io_enq_bits_opcode;
  wire [1:0] AsyncQueueSource_io_enq_bits_param;
  wire [1:0] AsyncQueueSource_io_enq_bits_size;
  wire  AsyncQueueSource_io_enq_bits_source;
  wire  AsyncQueueSource_io_enq_bits_sink;
  wire [31:0] AsyncQueueSource_io_enq_bits_data;
  wire  AsyncQueueSource_io_enq_bits_error;
  wire  AsyncQueueSource_io_ridx;
  wire  AsyncQueueSource_io_widx;
  wire [2:0] AsyncQueueSource_io_mem_0_opcode;
  wire [1:0] AsyncQueueSource_io_mem_0_param;
  wire [1:0] AsyncQueueSource_io_mem_0_size;
  wire  AsyncQueueSource_io_mem_0_source;
  wire  AsyncQueueSource_io_mem_0_sink;
  wire [31:0] AsyncQueueSource_io_mem_0_data;
  wire  AsyncQueueSource_io_mem_0_error;
  wire  AsyncQueueSource_io_sink_reset_n;
  wire  AsyncQueueSource_io_ridx_valid;
  wire  AsyncQueueSource_io_widx_valid;
  wire [2:0] _T_119_mem_0_opcode;
  wire [1:0] _T_119_mem_0_param;
  wire [1:0] _T_119_mem_0_size;
  wire  _T_119_mem_0_source;
  wire  _T_119_mem_0_sink;
  wire [31:0] _T_119_mem_0_data;
  wire  _T_119_mem_0_error;
  wire  _T_119_widx;
  wire  _T_119_widx_valid;
  wire  _T_125;
  AsyncQueueSink_1 AsyncQueueSink (
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits_opcode(AsyncQueueSink_io_deq_bits_opcode),
    .io_deq_bits_size(AsyncQueueSink_io_deq_bits_size),
    .io_deq_bits_source(AsyncQueueSink_io_deq_bits_source),
    .io_deq_bits_address(AsyncQueueSink_io_deq_bits_address),
    .io_deq_bits_mask(AsyncQueueSink_io_deq_bits_mask),
    .io_deq_bits_data(AsyncQueueSink_io_deq_bits_data),
    .io_ridx(AsyncQueueSink_io_ridx),
    .io_widx(AsyncQueueSink_io_widx),
    .io_mem_0_opcode(AsyncQueueSink_io_mem_0_opcode),
    .io_mem_0_size(AsyncQueueSink_io_mem_0_size),
    .io_mem_0_source(AsyncQueueSink_io_mem_0_source),
    .io_mem_0_address(AsyncQueueSink_io_mem_0_address),
    .io_mem_0_mask(AsyncQueueSink_io_mem_0_mask),
    .io_mem_0_data(AsyncQueueSink_io_mem_0_data),
    .io_source_reset_n(AsyncQueueSink_io_source_reset_n),
    .io_ridx_valid(AsyncQueueSink_io_ridx_valid),
    .io_widx_valid(AsyncQueueSink_io_widx_valid)
  );
  AsyncQueueSource_2 AsyncQueueSource (
    .clock(AsyncQueueSource_clock),
    .reset(AsyncQueueSource_reset),
    .io_enq_ready(AsyncQueueSource_io_enq_ready),
    .io_enq_valid(AsyncQueueSource_io_enq_valid),
    .io_enq_bits_opcode(AsyncQueueSource_io_enq_bits_opcode),
    .io_enq_bits_param(AsyncQueueSource_io_enq_bits_param),
    .io_enq_bits_size(AsyncQueueSource_io_enq_bits_size),
    .io_enq_bits_source(AsyncQueueSource_io_enq_bits_source),
    .io_enq_bits_sink(AsyncQueueSource_io_enq_bits_sink),
    .io_enq_bits_data(AsyncQueueSource_io_enq_bits_data),
    .io_enq_bits_error(AsyncQueueSource_io_enq_bits_error),
    .io_ridx(AsyncQueueSource_io_ridx),
    .io_widx(AsyncQueueSource_io_widx),
    .io_mem_0_opcode(AsyncQueueSource_io_mem_0_opcode),
    .io_mem_0_param(AsyncQueueSource_io_mem_0_param),
    .io_mem_0_size(AsyncQueueSource_io_mem_0_size),
    .io_mem_0_source(AsyncQueueSource_io_mem_0_source),
    .io_mem_0_sink(AsyncQueueSource_io_mem_0_sink),
    .io_mem_0_data(AsyncQueueSource_io_mem_0_data),
    .io_mem_0_error(AsyncQueueSource_io_mem_0_error),
    .io_sink_reset_n(AsyncQueueSource_io_sink_reset_n),
    .io_ridx_valid(AsyncQueueSource_io_ridx_valid),
    .io_widx_valid(AsyncQueueSource_io_widx_valid)
  );
  assign io_in_0_a_ridx = AsyncQueueSink_io_ridx;
  assign io_in_0_a_ridx_valid = AsyncQueueSink_io_ridx_valid;
  assign io_in_0_a_sink_reset_n = _T_105;
  assign io_in_0_d_mem_0_opcode = _T_119_mem_0_opcode;
  assign io_in_0_d_mem_0_param = _T_119_mem_0_param;
  assign io_in_0_d_mem_0_size = _T_119_mem_0_size;
  assign io_in_0_d_mem_0_source = _T_119_mem_0_source;
  assign io_in_0_d_mem_0_sink = _T_119_mem_0_sink;
  assign io_in_0_d_mem_0_data = _T_119_mem_0_data;
  assign io_in_0_d_mem_0_error = _T_119_mem_0_error;
  assign io_in_0_d_widx = _T_119_widx;
  assign io_in_0_d_widx_valid = _T_119_widx_valid;
  assign io_in_0_d_source_reset_n = _T_125;
  assign io_out_0_a_valid = _T_110_valid;
  assign io_out_0_a_bits_opcode = _T_110_bits_opcode;
  assign io_out_0_a_bits_size = _T_110_bits_size;
  assign io_out_0_a_bits_source = _T_110_bits_source;
  assign io_out_0_a_bits_address = _T_110_bits_address;
  assign io_out_0_a_bits_mask = _T_110_bits_mask;
  assign io_out_0_a_bits_data = _T_110_bits_data;
  assign io_out_0_d_ready = AsyncQueueSource_io_enq_ready;
  assign AsyncQueueSink_clock = clock;
  assign AsyncQueueSink_reset = reset;
  assign AsyncQueueSink_io_deq_ready = io_out_0_a_ready;
  assign AsyncQueueSink_io_widx = io_in_0_a_widx;
  assign AsyncQueueSink_io_mem_0_opcode = io_in_0_a_mem_0_opcode;
  assign AsyncQueueSink_io_mem_0_size = io_in_0_a_mem_0_size;
  assign AsyncQueueSink_io_mem_0_source = io_in_0_a_mem_0_source;
  assign AsyncQueueSink_io_mem_0_address = io_in_0_a_mem_0_address;
  assign AsyncQueueSink_io_mem_0_mask = io_in_0_a_mem_0_mask;
  assign AsyncQueueSink_io_mem_0_data = io_in_0_a_mem_0_data;
  assign AsyncQueueSink_io_source_reset_n = io_in_0_a_source_reset_n;
  assign AsyncQueueSink_io_widx_valid = io_in_0_a_widx_valid;
  assign _T_105 = AsyncQueueSink_reset == 1'h0;
  assign _T_110_valid = AsyncQueueSink_io_deq_valid;
  assign _T_110_bits_opcode = AsyncQueueSink_io_deq_bits_opcode;
  assign _T_110_bits_size = AsyncQueueSink_io_deq_bits_size;
  assign _T_110_bits_source = AsyncQueueSink_io_deq_bits_source;
  assign _T_110_bits_address = AsyncQueueSink_io_deq_bits_address;
  assign _T_110_bits_mask = AsyncQueueSink_io_deq_bits_mask;
  assign _T_110_bits_data = AsyncQueueSink_io_deq_bits_data;
  assign AsyncQueueSource_clock = clock;
  assign AsyncQueueSource_reset = reset;
  assign AsyncQueueSource_io_enq_valid = io_out_0_d_valid;
  assign AsyncQueueSource_io_enq_bits_opcode = io_out_0_d_bits_opcode;
  assign AsyncQueueSource_io_enq_bits_param = io_out_0_d_bits_param;
  assign AsyncQueueSource_io_enq_bits_size = io_out_0_d_bits_size;
  assign AsyncQueueSource_io_enq_bits_source = io_out_0_d_bits_source;
  assign AsyncQueueSource_io_enq_bits_sink = io_out_0_d_bits_sink;
  assign AsyncQueueSource_io_enq_bits_data = io_out_0_d_bits_data;
  assign AsyncQueueSource_io_enq_bits_error = io_out_0_d_bits_error;
  assign AsyncQueueSource_io_ridx = io_in_0_d_ridx;
  assign AsyncQueueSource_io_sink_reset_n = io_in_0_d_sink_reset_n;
  assign AsyncQueueSource_io_ridx_valid = io_in_0_d_ridx_valid;
  assign _T_119_mem_0_opcode = AsyncQueueSource_io_mem_0_opcode;
  assign _T_119_mem_0_param = AsyncQueueSource_io_mem_0_param;
  assign _T_119_mem_0_size = AsyncQueueSource_io_mem_0_size;
  assign _T_119_mem_0_source = AsyncQueueSource_io_mem_0_source;
  assign _T_119_mem_0_sink = AsyncQueueSource_io_mem_0_sink;
  assign _T_119_mem_0_data = AsyncQueueSource_io_mem_0_data;
  assign _T_119_mem_0_error = AsyncQueueSource_io_mem_0_error;
  assign _T_119_widx = AsyncQueueSource_io_widx;
  assign _T_119_widx_valid = AsyncQueueSource_io_widx_valid;
  assign _T_125 = AsyncQueueSource_reset == 1'h0;
endmodule
module AsyncQueueSink_2(
  input        clock,
  input        reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output       io_deq_bits_resumereq,
  output [9:0] io_deq_bits_hartsel,
  output       io_ridx,
  input        io_widx,
  input        io_mem_0_resumereq,
  input  [9:0] io_mem_0_hartsel,
  input        io_source_reset_n,
  output       io_ridx_valid,
  input        io_widx_valid
);
  wire  source_ready;
  wire  _T_17;
  wire  _T_19;
  wire  ridx_bin_clock;
  wire  ridx_bin_reset;
  wire  ridx_bin_io_d;
  wire  ridx_bin_io_q;
  wire  ridx_bin_io_en;
  wire [1:0] _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_28;
  wire  ridx;
  wire  widx_gray_sync_0_clock;
  wire  widx_gray_sync_0_reset;
  wire  widx_gray_sync_0_io_d;
  wire  widx_gray_sync_0_io_q;
  wire  widx_gray_sync_0_io_en;
  wire  widx_gray_sync_1_clock;
  wire  widx_gray_sync_1_reset;
  wire  widx_gray_sync_1_io_d;
  wire  widx_gray_sync_1_io_q;
  wire  widx_gray_sync_1_io_en;
  wire  widx_gray_sync_2_clock;
  wire  widx_gray_sync_2_reset;
  wire  widx_gray_sync_2_io_d;
  wire  widx_gray_sync_2_io_q;
  wire  widx_gray_sync_2_io_en;
  wire  _T_32;
  wire  valid;
  reg  _T_36_resumereq;
  reg [31:0] _RAND_0;
  reg [9:0] _T_36_hartsel;
  reg [31:0] _RAND_1;
  wire  _GEN_0;
  wire [9:0] _GEN_1;
  wire  valid_reg_clock;
  wire  valid_reg_reset;
  wire  valid_reg_io_d;
  wire  valid_reg_io_q;
  wire  valid_reg_io_en;
  wire  valid_reg_1;
  wire  _T_38;
  wire  ridx_gray_clock;
  wire  ridx_gray_reset;
  wire  ridx_gray_io_d;
  wire  ridx_gray_io_q;
  wire  ridx_gray_io_en;
  wire  AsyncValidSync_clock;
  wire  AsyncValidSync_reset;
  wire  AsyncValidSync_io_in;
  wire  AsyncValidSync_io_out;
  wire  AsyncValidSync_1_clock;
  wire  AsyncValidSync_1_reset;
  wire  AsyncValidSync_1_io_in;
  wire  AsyncValidSync_1_io_out;
  wire  AsyncValidSync_2_clock;
  wire  AsyncValidSync_2_reset;
  wire  AsyncValidSync_2_io_in;
  wire  AsyncValidSync_2_io_out;
  wire  _T_42;
  wire  _T_43;
  wire  _T_60;
  wire  AsyncResetRegVec_clock;
  wire  AsyncResetRegVec_reset;
  wire  AsyncResetRegVec_io_d;
  wire  AsyncResetRegVec_io_q;
  wire  AsyncResetRegVec_io_en;
  AsyncResetRegVec_1 ridx_bin (
    .clock(ridx_bin_clock),
    .reset(ridx_bin_reset),
    .io_d(ridx_bin_io_d),
    .io_q(ridx_bin_io_q),
    .io_en(ridx_bin_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_0 (
    .clock(widx_gray_sync_0_clock),
    .reset(widx_gray_sync_0_reset),
    .io_d(widx_gray_sync_0_io_d),
    .io_q(widx_gray_sync_0_io_q),
    .io_en(widx_gray_sync_0_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_1 (
    .clock(widx_gray_sync_1_clock),
    .reset(widx_gray_sync_1_reset),
    .io_d(widx_gray_sync_1_io_d),
    .io_q(widx_gray_sync_1_io_q),
    .io_en(widx_gray_sync_1_io_en)
  );
  AsyncResetRegVec_1 widx_gray_sync_2 (
    .clock(widx_gray_sync_2_clock),
    .reset(widx_gray_sync_2_reset),
    .io_d(widx_gray_sync_2_io_d),
    .io_q(widx_gray_sync_2_io_q),
    .io_en(widx_gray_sync_2_io_en)
  );
  AsyncResetRegVec_1 valid_reg (
    .clock(valid_reg_clock),
    .reset(valid_reg_reset),
    .io_d(valid_reg_io_d),
    .io_q(valid_reg_io_q),
    .io_en(valid_reg_io_en)
  );
  AsyncResetRegVec_1 ridx_gray (
    .clock(ridx_gray_clock),
    .reset(ridx_gray_reset),
    .io_d(ridx_gray_io_d),
    .io_q(ridx_gray_io_q),
    .io_en(ridx_gray_io_en)
  );
  AsyncValidSync_3 AsyncValidSync (
    .clock(AsyncValidSync_clock),
    .reset(AsyncValidSync_reset),
    .io_in(AsyncValidSync_io_in),
    .io_out(AsyncValidSync_io_out)
  );
  AsyncValidSync_4 AsyncValidSync_1 (
    .clock(AsyncValidSync_1_clock),
    .reset(AsyncValidSync_1_reset),
    .io_in(AsyncValidSync_1_io_in),
    .io_out(AsyncValidSync_1_io_out)
  );
  AsyncValidSync_5 AsyncValidSync_2 (
    .clock(AsyncValidSync_2_clock),
    .reset(AsyncValidSync_2_reset),
    .io_in(AsyncValidSync_2_io_in),
    .io_out(AsyncValidSync_2_io_out)
  );
  AsyncResetRegVec_1 AsyncResetRegVec (
    .clock(AsyncResetRegVec_clock),
    .reset(AsyncResetRegVec_reset),
    .io_d(AsyncResetRegVec_io_d),
    .io_q(AsyncResetRegVec_io_q),
    .io_en(AsyncResetRegVec_io_en)
  );
  assign io_deq_valid = _T_38;
  assign io_deq_bits_resumereq = _T_36_resumereq;
  assign io_deq_bits_hartsel = _T_36_hartsel;
  assign io_ridx = ridx_gray_io_q;
  assign io_ridx_valid = AsyncValidSync_io_out;
  assign source_ready = AsyncValidSync_2_io_out;
  assign _T_17 = io_deq_ready & io_deq_valid;
  assign _T_19 = source_ready == 1'h0;
  assign ridx_bin_clock = clock;
  assign ridx_bin_reset = reset;
  assign ridx_bin_io_d = _T_26;
  assign ridx_bin_io_en = 1'h1;
  assign _T_24 = ridx_bin_io_q + _T_17;
  assign _T_25 = _T_24[0:0];
  assign _T_26 = _T_19 ? 1'h0 : _T_25;
  assign _T_28 = _T_26 >> 1'h1;
  assign ridx = _T_26 ^ _T_28;
  assign widx_gray_sync_0_clock = clock;
  assign widx_gray_sync_0_reset = reset;
  assign widx_gray_sync_0_io_d = widx_gray_sync_1_io_q;
  assign widx_gray_sync_0_io_en = 1'h1;
  assign widx_gray_sync_1_clock = clock;
  assign widx_gray_sync_1_reset = reset;
  assign widx_gray_sync_1_io_d = widx_gray_sync_2_io_q;
  assign widx_gray_sync_1_io_en = 1'h1;
  assign widx_gray_sync_2_clock = clock;
  assign widx_gray_sync_2_reset = reset;
  assign widx_gray_sync_2_io_d = io_widx;
  assign widx_gray_sync_2_io_en = 1'h1;
  assign _T_32 = ridx != widx_gray_sync_0_io_q;
  assign valid = source_ready & _T_32;
  assign _GEN_0 = valid ? io_mem_0_resumereq : _T_36_resumereq;
  assign _GEN_1 = valid ? io_mem_0_hartsel : _T_36_hartsel;
  assign valid_reg_clock = clock;
  assign valid_reg_reset = reset;
  assign valid_reg_io_d = valid;
  assign valid_reg_io_en = 1'h1;
  assign valid_reg_1 = valid_reg_io_q;
  assign _T_38 = valid_reg_1 & source_ready;
  assign ridx_gray_clock = clock;
  assign ridx_gray_reset = reset;
  assign ridx_gray_io_d = ridx;
  assign ridx_gray_io_en = 1'h1;
  assign AsyncValidSync_clock = clock;
  assign AsyncValidSync_reset = _T_43;
  assign AsyncValidSync_io_in = 1'h1;
  assign AsyncValidSync_1_clock = clock;
  assign AsyncValidSync_1_reset = _T_43;
  assign AsyncValidSync_1_io_in = io_widx_valid;
  assign AsyncValidSync_2_clock = clock;
  assign AsyncValidSync_2_reset = reset;
  assign AsyncValidSync_2_io_in = AsyncValidSync_1_io_out;
  assign _T_42 = io_source_reset_n == 1'h0;
  assign _T_43 = reset | _T_42;
  assign _T_60 = io_widx == io_ridx;
  assign AsyncResetRegVec_clock = clock;
  assign AsyncResetRegVec_reset = reset;
  assign AsyncResetRegVec_io_d = _T_60;
  assign AsyncResetRegVec_io_en = 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_36_resumereq = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_36_hartsel = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (valid) begin
      _T_36_resumereq <= io_mem_0_resumereq;
    end
    if (valid) begin
      _T_36_hartsel <= io_mem_0_hartsel;
    end
  end
endmodule
module AsyncResetRegVec_89(
  input        clock,
  input        reset,
  input  [2:0] io_d,
  output [2:0] io_q,
  input        io_en
);
  wire  reg_0_rst;
  wire  reg_0_clk;
  wire  reg_0_en;
  wire  reg_0_q;
  wire  reg_0_d;
  wire  reg_1_rst;
  wire  reg_1_clk;
  wire  reg_1_en;
  wire  reg_1_q;
  wire  reg_1_d;
  wire  reg_2_rst;
  wire  reg_2_clk;
  wire  reg_2_en;
  wire  reg_2_q;
  wire  reg_2_d;
  wire  _T_5;
  wire  _T_6;
  wire  _T_7;
  wire [1:0] _T_8;
  wire [2:0] _T_9;
  AsyncResetReg reg_0 (
    .rst(reg_0_rst),
    .clk(reg_0_clk),
    .en(reg_0_en),
    .q(reg_0_q),
    .d(reg_0_d)
  );
  AsyncResetReg reg_1 (
    .rst(reg_1_rst),
    .clk(reg_1_clk),
    .en(reg_1_en),
    .q(reg_1_q),
    .d(reg_1_d)
  );
  AsyncResetReg reg_2 (
    .rst(reg_2_rst),
    .clk(reg_2_clk),
    .en(reg_2_en),
    .q(reg_2_q),
    .d(reg_2_d)
  );
  assign io_q = _T_9;
  assign reg_0_rst = reset;
  assign reg_0_clk = clock;
  assign reg_0_en = io_en;
  assign reg_0_d = _T_5;
  assign reg_1_rst = reset;
  assign reg_1_clk = clock;
  assign reg_1_en = io_en;
  assign reg_1_d = _T_6;
  assign reg_2_rst = reset;
  assign reg_2_clk = clock;
  assign reg_2_en = io_en;
  assign reg_2_d = _T_7;
  assign _T_5 = io_d[0];
  assign _T_6 = io_d[1];
  assign _T_7 = io_d[2];
  assign _T_8 = {reg_2_q,reg_1_q};
  assign _T_9 = {_T_8,reg_0_q};
endmodule
module ResetCatchAndSync(
  input   clock,
  input   reset,
  output  io_sync_reset
);
  wire  reset_n_catch_reg_clock;
  wire  reset_n_catch_reg_reset;
  wire [2:0] reset_n_catch_reg_io_d;
  wire [2:0] reset_n_catch_reg_io_q;
  wire  reset_n_catch_reg_io_en;
  wire [1:0] _T_5;
  wire [2:0] _T_6;
  wire  _T_7;
  wire  _T_8;
  AsyncResetRegVec_89 reset_n_catch_reg (
    .clock(reset_n_catch_reg_clock),
    .reset(reset_n_catch_reg_reset),
    .io_d(reset_n_catch_reg_io_d),
    .io_q(reset_n_catch_reg_io_q),
    .io_en(reset_n_catch_reg_io_en)
  );
  assign io_sync_reset = _T_8;
  assign reset_n_catch_reg_clock = clock;
  assign reset_n_catch_reg_reset = reset;
  assign reset_n_catch_reg_io_d = _T_6;
  assign reset_n_catch_reg_io_en = 1'h1;
  assign _T_5 = reset_n_catch_reg_io_q[2:1];
  assign _T_6 = {1'h1,_T_5};
  assign _T_7 = reset_n_catch_reg_io_q[0];
  assign _T_8 = ~ _T_7;
endmodule
module TLDebugModuleInnerAsync_dmInner(
  input         clock,
  input         reset,
  input  [2:0]  io_dmi_in_0_a_mem_0_opcode,
  input  [1:0]  io_dmi_in_0_a_mem_0_size,
  input         io_dmi_in_0_a_mem_0_source,
  input  [8:0]  io_dmi_in_0_a_mem_0_address,
  input  [3:0]  io_dmi_in_0_a_mem_0_mask,
  input  [31:0] io_dmi_in_0_a_mem_0_data,
  output        io_dmi_in_0_a_ridx,
  input         io_dmi_in_0_a_widx,
  output        io_dmi_in_0_a_ridx_valid,
  input         io_dmi_in_0_a_widx_valid,
  input         io_dmi_in_0_a_source_reset_n,
  output        io_dmi_in_0_a_sink_reset_n,
  output [2:0]  io_dmi_in_0_d_mem_0_opcode,
  output [1:0]  io_dmi_in_0_d_mem_0_param,
  output [1:0]  io_dmi_in_0_d_mem_0_size,
  output        io_dmi_in_0_d_mem_0_source,
  output        io_dmi_in_0_d_mem_0_sink,
  output [31:0] io_dmi_in_0_d_mem_0_data,
  output        io_dmi_in_0_d_mem_0_error,
  input         io_dmi_in_0_d_ridx,
  output        io_dmi_in_0_d_widx,
  input         io_dmi_in_0_d_ridx_valid,
  output        io_dmi_in_0_d_widx_valid,
  output        io_dmi_in_0_d_source_reset_n,
  input         io_dmi_in_0_d_sink_reset_n,
  output        io_tl_in_0_a_ready,
  input         io_tl_in_0_a_valid,
  input  [2:0]  io_tl_in_0_a_bits_opcode,
  input  [1:0]  io_tl_in_0_a_bits_size,
  input  [9:0]  io_tl_in_0_a_bits_source,
  input  [11:0] io_tl_in_0_a_bits_address,
  input  [3:0]  io_tl_in_0_a_bits_mask,
  input  [31:0] io_tl_in_0_a_bits_data,
  input         io_tl_in_0_d_ready,
  output        io_tl_in_0_d_valid,
  output [2:0]  io_tl_in_0_d_bits_opcode,
  output [1:0]  io_tl_in_0_d_bits_param,
  output [1:0]  io_tl_in_0_d_bits_size,
  output [9:0]  io_tl_in_0_d_bits_source,
  output        io_tl_in_0_d_bits_sink,
  output [31:0] io_tl_in_0_d_bits_data,
  output        io_tl_in_0_d_bits_error,
  input         io_dmactive,
  input         io_innerCtrl_mem_0_resumereq,
  input  [9:0]  io_innerCtrl_mem_0_hartsel,
  output        io_innerCtrl_ridx,
  input         io_innerCtrl_widx,
  output        io_innerCtrl_ridx_valid,
  input         io_innerCtrl_widx_valid,
  input         io_innerCtrl_source_reset_n,
  output        io_innerCtrl_sink_reset_n,
  input         io_debugUnavail_0
);
  wire  dmInner_clock;
  wire  dmInner_reset;
  wire  dmInner_io_hart_in_0_a_ready;
  wire  dmInner_io_hart_in_0_a_valid;
  wire [2:0] dmInner_io_hart_in_0_a_bits_opcode;
  wire [1:0] dmInner_io_hart_in_0_a_bits_size;
  wire [9:0] dmInner_io_hart_in_0_a_bits_source;
  wire [11:0] dmInner_io_hart_in_0_a_bits_address;
  wire [3:0] dmInner_io_hart_in_0_a_bits_mask;
  wire [31:0] dmInner_io_hart_in_0_a_bits_data;
  wire  dmInner_io_hart_in_0_d_ready;
  wire  dmInner_io_hart_in_0_d_valid;
  wire [2:0] dmInner_io_hart_in_0_d_bits_opcode;
  wire [1:0] dmInner_io_hart_in_0_d_bits_param;
  wire [1:0] dmInner_io_hart_in_0_d_bits_size;
  wire [9:0] dmInner_io_hart_in_0_d_bits_source;
  wire  dmInner_io_hart_in_0_d_bits_sink;
  wire [31:0] dmInner_io_hart_in_0_d_bits_data;
  wire  dmInner_io_hart_in_0_d_bits_error;
  wire  dmInner_io_dmi_in_0_a_ready;
  wire  dmInner_io_dmi_in_0_a_valid;
  wire [2:0] dmInner_io_dmi_in_0_a_bits_opcode;
  wire [1:0] dmInner_io_dmi_in_0_a_bits_size;
  wire  dmInner_io_dmi_in_0_a_bits_source;
  wire [8:0] dmInner_io_dmi_in_0_a_bits_address;
  wire [3:0] dmInner_io_dmi_in_0_a_bits_mask;
  wire [31:0] dmInner_io_dmi_in_0_a_bits_data;
  wire  dmInner_io_dmi_in_0_d_ready;
  wire  dmInner_io_dmi_in_0_d_valid;
  wire [2:0] dmInner_io_dmi_in_0_d_bits_opcode;
  wire [1:0] dmInner_io_dmi_in_0_d_bits_param;
  wire [1:0] dmInner_io_dmi_in_0_d_bits_size;
  wire  dmInner_io_dmi_in_0_d_bits_source;
  wire  dmInner_io_dmi_in_0_d_bits_sink;
  wire [31:0] dmInner_io_dmi_in_0_d_bits_data;
  wire  dmInner_io_dmi_in_0_d_bits_error;
  wire  dmInner_io_dmactive;
  wire  dmInner_io_innerCtrl_ready;
  wire  dmInner_io_innerCtrl_valid;
  wire  dmInner_io_innerCtrl_bits_resumereq;
  wire [9:0] dmInner_io_innerCtrl_bits_hartsel;
  wire  dmInner_io_debugUnavail_0;
  wire  TLAsyncCrossingSink_clock;
  wire  TLAsyncCrossingSink_reset;
  wire [2:0] TLAsyncCrossingSink_io_in_0_a_mem_0_opcode;
  wire [1:0] TLAsyncCrossingSink_io_in_0_a_mem_0_size;
  wire  TLAsyncCrossingSink_io_in_0_a_mem_0_source;
  wire [8:0] TLAsyncCrossingSink_io_in_0_a_mem_0_address;
  wire [3:0] TLAsyncCrossingSink_io_in_0_a_mem_0_mask;
  wire [31:0] TLAsyncCrossingSink_io_in_0_a_mem_0_data;
  wire  TLAsyncCrossingSink_io_in_0_a_ridx;
  wire  TLAsyncCrossingSink_io_in_0_a_widx;
  wire  TLAsyncCrossingSink_io_in_0_a_ridx_valid;
  wire  TLAsyncCrossingSink_io_in_0_a_widx_valid;
  wire  TLAsyncCrossingSink_io_in_0_a_source_reset_n;
  wire  TLAsyncCrossingSink_io_in_0_a_sink_reset_n;
  wire [2:0] TLAsyncCrossingSink_io_in_0_d_mem_0_opcode;
  wire [1:0] TLAsyncCrossingSink_io_in_0_d_mem_0_param;
  wire [1:0] TLAsyncCrossingSink_io_in_0_d_mem_0_size;
  wire  TLAsyncCrossingSink_io_in_0_d_mem_0_source;
  wire  TLAsyncCrossingSink_io_in_0_d_mem_0_sink;
  wire [31:0] TLAsyncCrossingSink_io_in_0_d_mem_0_data;
  wire  TLAsyncCrossingSink_io_in_0_d_mem_0_error;
  wire  TLAsyncCrossingSink_io_in_0_d_ridx;
  wire  TLAsyncCrossingSink_io_in_0_d_widx;
  wire  TLAsyncCrossingSink_io_in_0_d_ridx_valid;
  wire  TLAsyncCrossingSink_io_in_0_d_widx_valid;
  wire  TLAsyncCrossingSink_io_in_0_d_source_reset_n;
  wire  TLAsyncCrossingSink_io_in_0_d_sink_reset_n;
  wire  TLAsyncCrossingSink_io_out_0_a_ready;
  wire  TLAsyncCrossingSink_io_out_0_a_valid;
  wire [2:0] TLAsyncCrossingSink_io_out_0_a_bits_opcode;
  wire [1:0] TLAsyncCrossingSink_io_out_0_a_bits_size;
  wire  TLAsyncCrossingSink_io_out_0_a_bits_source;
  wire [8:0] TLAsyncCrossingSink_io_out_0_a_bits_address;
  wire [3:0] TLAsyncCrossingSink_io_out_0_a_bits_mask;
  wire [31:0] TLAsyncCrossingSink_io_out_0_a_bits_data;
  wire  TLAsyncCrossingSink_io_out_0_d_ready;
  wire  TLAsyncCrossingSink_io_out_0_d_valid;
  wire [2:0] TLAsyncCrossingSink_io_out_0_d_bits_opcode;
  wire [1:0] TLAsyncCrossingSink_io_out_0_d_bits_param;
  wire [1:0] TLAsyncCrossingSink_io_out_0_d_bits_size;
  wire  TLAsyncCrossingSink_io_out_0_d_bits_source;
  wire  TLAsyncCrossingSink_io_out_0_d_bits_sink;
  wire [31:0] TLAsyncCrossingSink_io_out_0_d_bits_data;
  wire  TLAsyncCrossingSink_io_out_0_d_bits_error;
  wire  AsyncQueueSink_clock;
  wire  AsyncQueueSink_reset;
  wire  AsyncQueueSink_io_deq_ready;
  wire  AsyncQueueSink_io_deq_valid;
  wire  AsyncQueueSink_io_deq_bits_resumereq;
  wire [9:0] AsyncQueueSink_io_deq_bits_hartsel;
  wire  AsyncQueueSink_io_ridx;
  wire  AsyncQueueSink_io_widx;
  wire  AsyncQueueSink_io_mem_0_resumereq;
  wire [9:0] AsyncQueueSink_io_mem_0_hartsel;
  wire  AsyncQueueSink_io_source_reset_n;
  wire  AsyncQueueSink_io_ridx_valid;
  wire  AsyncQueueSink_io_widx_valid;
  wire  _T_154;
  wire  _T_159_ready;
  wire  _T_159_valid;
  wire  _T_159_bits_resumereq;
  wire [9:0] _T_159_bits_hartsel;
  wire  _T_163;
  wire  ResetCatchAndSync_clock;
  wire  ResetCatchAndSync_reset;
  wire  ResetCatchAndSync_io_sync_reset;
  wire  _T_164;
  TLDebugModuleInner_dmInner dmInner (
    .clock(dmInner_clock),
    .reset(dmInner_reset),
    .io_hart_in_0_a_ready(dmInner_io_hart_in_0_a_ready),
    .io_hart_in_0_a_valid(dmInner_io_hart_in_0_a_valid),
    .io_hart_in_0_a_bits_opcode(dmInner_io_hart_in_0_a_bits_opcode),
    .io_hart_in_0_a_bits_size(dmInner_io_hart_in_0_a_bits_size),
    .io_hart_in_0_a_bits_source(dmInner_io_hart_in_0_a_bits_source),
    .io_hart_in_0_a_bits_address(dmInner_io_hart_in_0_a_bits_address),
    .io_hart_in_0_a_bits_mask(dmInner_io_hart_in_0_a_bits_mask),
    .io_hart_in_0_a_bits_data(dmInner_io_hart_in_0_a_bits_data),
    .io_hart_in_0_d_ready(dmInner_io_hart_in_0_d_ready),
    .io_hart_in_0_d_valid(dmInner_io_hart_in_0_d_valid),
    .io_hart_in_0_d_bits_opcode(dmInner_io_hart_in_0_d_bits_opcode),
    .io_hart_in_0_d_bits_param(dmInner_io_hart_in_0_d_bits_param),
    .io_hart_in_0_d_bits_size(dmInner_io_hart_in_0_d_bits_size),
    .io_hart_in_0_d_bits_source(dmInner_io_hart_in_0_d_bits_source),
    .io_hart_in_0_d_bits_sink(dmInner_io_hart_in_0_d_bits_sink),
    .io_hart_in_0_d_bits_data(dmInner_io_hart_in_0_d_bits_data),
    .io_hart_in_0_d_bits_error(dmInner_io_hart_in_0_d_bits_error),
    .io_dmi_in_0_a_ready(dmInner_io_dmi_in_0_a_ready),
    .io_dmi_in_0_a_valid(dmInner_io_dmi_in_0_a_valid),
    .io_dmi_in_0_a_bits_opcode(dmInner_io_dmi_in_0_a_bits_opcode),
    .io_dmi_in_0_a_bits_size(dmInner_io_dmi_in_0_a_bits_size),
    .io_dmi_in_0_a_bits_source(dmInner_io_dmi_in_0_a_bits_source),
    .io_dmi_in_0_a_bits_address(dmInner_io_dmi_in_0_a_bits_address),
    .io_dmi_in_0_a_bits_mask(dmInner_io_dmi_in_0_a_bits_mask),
    .io_dmi_in_0_a_bits_data(dmInner_io_dmi_in_0_a_bits_data),
    .io_dmi_in_0_d_ready(dmInner_io_dmi_in_0_d_ready),
    .io_dmi_in_0_d_valid(dmInner_io_dmi_in_0_d_valid),
    .io_dmi_in_0_d_bits_opcode(dmInner_io_dmi_in_0_d_bits_opcode),
    .io_dmi_in_0_d_bits_param(dmInner_io_dmi_in_0_d_bits_param),
    .io_dmi_in_0_d_bits_size(dmInner_io_dmi_in_0_d_bits_size),
    .io_dmi_in_0_d_bits_source(dmInner_io_dmi_in_0_d_bits_source),
    .io_dmi_in_0_d_bits_sink(dmInner_io_dmi_in_0_d_bits_sink),
    .io_dmi_in_0_d_bits_data(dmInner_io_dmi_in_0_d_bits_data),
    .io_dmi_in_0_d_bits_error(dmInner_io_dmi_in_0_d_bits_error),
    .io_dmactive(dmInner_io_dmactive),
    .io_innerCtrl_ready(dmInner_io_innerCtrl_ready),
    .io_innerCtrl_valid(dmInner_io_innerCtrl_valid),
    .io_innerCtrl_bits_resumereq(dmInner_io_innerCtrl_bits_resumereq),
    .io_innerCtrl_bits_hartsel(dmInner_io_innerCtrl_bits_hartsel),
    .io_debugUnavail_0(dmInner_io_debugUnavail_0)
  );
  TLAsyncCrossingSink TLAsyncCrossingSink (
    .clock(TLAsyncCrossingSink_clock),
    .reset(TLAsyncCrossingSink_reset),
    .io_in_0_a_mem_0_opcode(TLAsyncCrossingSink_io_in_0_a_mem_0_opcode),
    .io_in_0_a_mem_0_size(TLAsyncCrossingSink_io_in_0_a_mem_0_size),
    .io_in_0_a_mem_0_source(TLAsyncCrossingSink_io_in_0_a_mem_0_source),
    .io_in_0_a_mem_0_address(TLAsyncCrossingSink_io_in_0_a_mem_0_address),
    .io_in_0_a_mem_0_mask(TLAsyncCrossingSink_io_in_0_a_mem_0_mask),
    .io_in_0_a_mem_0_data(TLAsyncCrossingSink_io_in_0_a_mem_0_data),
    .io_in_0_a_ridx(TLAsyncCrossingSink_io_in_0_a_ridx),
    .io_in_0_a_widx(TLAsyncCrossingSink_io_in_0_a_widx),
    .io_in_0_a_ridx_valid(TLAsyncCrossingSink_io_in_0_a_ridx_valid),
    .io_in_0_a_widx_valid(TLAsyncCrossingSink_io_in_0_a_widx_valid),
    .io_in_0_a_source_reset_n(TLAsyncCrossingSink_io_in_0_a_source_reset_n),
    .io_in_0_a_sink_reset_n(TLAsyncCrossingSink_io_in_0_a_sink_reset_n),
    .io_in_0_d_mem_0_opcode(TLAsyncCrossingSink_io_in_0_d_mem_0_opcode),
    .io_in_0_d_mem_0_param(TLAsyncCrossingSink_io_in_0_d_mem_0_param),
    .io_in_0_d_mem_0_size(TLAsyncCrossingSink_io_in_0_d_mem_0_size),
    .io_in_0_d_mem_0_source(TLAsyncCrossingSink_io_in_0_d_mem_0_source),
    .io_in_0_d_mem_0_sink(TLAsyncCrossingSink_io_in_0_d_mem_0_sink),
    .io_in_0_d_mem_0_data(TLAsyncCrossingSink_io_in_0_d_mem_0_data),
    .io_in_0_d_mem_0_error(TLAsyncCrossingSink_io_in_0_d_mem_0_error),
    .io_in_0_d_ridx(TLAsyncCrossingSink_io_in_0_d_ridx),
    .io_in_0_d_widx(TLAsyncCrossingSink_io_in_0_d_widx),
    .io_in_0_d_ridx_valid(TLAsyncCrossingSink_io_in_0_d_ridx_valid),
    .io_in_0_d_widx_valid(TLAsyncCrossingSink_io_in_0_d_widx_valid),
    .io_in_0_d_source_reset_n(TLAsyncCrossingSink_io_in_0_d_source_reset_n),
    .io_in_0_d_sink_reset_n(TLAsyncCrossingSink_io_in_0_d_sink_reset_n),
    .io_out_0_a_ready(TLAsyncCrossingSink_io_out_0_a_ready),
    .io_out_0_a_valid(TLAsyncCrossingSink_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLAsyncCrossingSink_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(TLAsyncCrossingSink_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLAsyncCrossingSink_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLAsyncCrossingSink_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLAsyncCrossingSink_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLAsyncCrossingSink_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLAsyncCrossingSink_io_out_0_d_ready),
    .io_out_0_d_valid(TLAsyncCrossingSink_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLAsyncCrossingSink_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLAsyncCrossingSink_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLAsyncCrossingSink_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLAsyncCrossingSink_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLAsyncCrossingSink_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLAsyncCrossingSink_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLAsyncCrossingSink_io_out_0_d_bits_error)
  );
  AsyncQueueSink_2 AsyncQueueSink (
    .clock(AsyncQueueSink_clock),
    .reset(AsyncQueueSink_reset),
    .io_deq_ready(AsyncQueueSink_io_deq_ready),
    .io_deq_valid(AsyncQueueSink_io_deq_valid),
    .io_deq_bits_resumereq(AsyncQueueSink_io_deq_bits_resumereq),
    .io_deq_bits_hartsel(AsyncQueueSink_io_deq_bits_hartsel),
    .io_ridx(AsyncQueueSink_io_ridx),
    .io_widx(AsyncQueueSink_io_widx),
    .io_mem_0_resumereq(AsyncQueueSink_io_mem_0_resumereq),
    .io_mem_0_hartsel(AsyncQueueSink_io_mem_0_hartsel),
    .io_source_reset_n(AsyncQueueSink_io_source_reset_n),
    .io_ridx_valid(AsyncQueueSink_io_ridx_valid),
    .io_widx_valid(AsyncQueueSink_io_widx_valid)
  );
  ResetCatchAndSync ResetCatchAndSync (
    .clock(ResetCatchAndSync_clock),
    .reset(ResetCatchAndSync_reset),
    .io_sync_reset(ResetCatchAndSync_io_sync_reset)
  );
  assign io_dmi_in_0_a_ridx = TLAsyncCrossingSink_io_in_0_a_ridx;
  assign io_dmi_in_0_a_ridx_valid = TLAsyncCrossingSink_io_in_0_a_ridx_valid;
  assign io_dmi_in_0_a_sink_reset_n = TLAsyncCrossingSink_io_in_0_a_sink_reset_n;
  assign io_dmi_in_0_d_mem_0_opcode = TLAsyncCrossingSink_io_in_0_d_mem_0_opcode;
  assign io_dmi_in_0_d_mem_0_param = TLAsyncCrossingSink_io_in_0_d_mem_0_param;
  assign io_dmi_in_0_d_mem_0_size = TLAsyncCrossingSink_io_in_0_d_mem_0_size;
  assign io_dmi_in_0_d_mem_0_source = TLAsyncCrossingSink_io_in_0_d_mem_0_source;
  assign io_dmi_in_0_d_mem_0_sink = TLAsyncCrossingSink_io_in_0_d_mem_0_sink;
  assign io_dmi_in_0_d_mem_0_data = TLAsyncCrossingSink_io_in_0_d_mem_0_data;
  assign io_dmi_in_0_d_mem_0_error = TLAsyncCrossingSink_io_in_0_d_mem_0_error;
  assign io_dmi_in_0_d_widx = TLAsyncCrossingSink_io_in_0_d_widx;
  assign io_dmi_in_0_d_widx_valid = TLAsyncCrossingSink_io_in_0_d_widx_valid;
  assign io_dmi_in_0_d_source_reset_n = TLAsyncCrossingSink_io_in_0_d_source_reset_n;
  assign io_tl_in_0_a_ready = dmInner_io_hart_in_0_a_ready;
  assign io_tl_in_0_d_valid = dmInner_io_hart_in_0_d_valid;
  assign io_tl_in_0_d_bits_opcode = dmInner_io_hart_in_0_d_bits_opcode;
  assign io_tl_in_0_d_bits_param = dmInner_io_hart_in_0_d_bits_param;
  assign io_tl_in_0_d_bits_size = dmInner_io_hart_in_0_d_bits_size;
  assign io_tl_in_0_d_bits_source = dmInner_io_hart_in_0_d_bits_source;
  assign io_tl_in_0_d_bits_sink = dmInner_io_hart_in_0_d_bits_sink;
  assign io_tl_in_0_d_bits_data = dmInner_io_hart_in_0_d_bits_data;
  assign io_tl_in_0_d_bits_error = dmInner_io_hart_in_0_d_bits_error;
  assign io_innerCtrl_ridx = AsyncQueueSink_io_ridx;
  assign io_innerCtrl_ridx_valid = AsyncQueueSink_io_ridx_valid;
  assign io_innerCtrl_sink_reset_n = _T_154;
  assign dmInner_clock = clock;
  assign dmInner_reset = reset;
  assign dmInner_io_hart_in_0_a_valid = io_tl_in_0_a_valid;
  assign dmInner_io_hart_in_0_a_bits_opcode = io_tl_in_0_a_bits_opcode;
  assign dmInner_io_hart_in_0_a_bits_size = io_tl_in_0_a_bits_size;
  assign dmInner_io_hart_in_0_a_bits_source = io_tl_in_0_a_bits_source;
  assign dmInner_io_hart_in_0_a_bits_address = io_tl_in_0_a_bits_address;
  assign dmInner_io_hart_in_0_a_bits_mask = io_tl_in_0_a_bits_mask;
  assign dmInner_io_hart_in_0_a_bits_data = io_tl_in_0_a_bits_data;
  assign dmInner_io_hart_in_0_d_ready = io_tl_in_0_d_ready;
  assign dmInner_io_dmi_in_0_a_valid = TLAsyncCrossingSink_io_out_0_a_valid;
  assign dmInner_io_dmi_in_0_a_bits_opcode = TLAsyncCrossingSink_io_out_0_a_bits_opcode;
  assign dmInner_io_dmi_in_0_a_bits_size = TLAsyncCrossingSink_io_out_0_a_bits_size;
  assign dmInner_io_dmi_in_0_a_bits_source = TLAsyncCrossingSink_io_out_0_a_bits_source;
  assign dmInner_io_dmi_in_0_a_bits_address = TLAsyncCrossingSink_io_out_0_a_bits_address;
  assign dmInner_io_dmi_in_0_a_bits_mask = TLAsyncCrossingSink_io_out_0_a_bits_mask;
  assign dmInner_io_dmi_in_0_a_bits_data = TLAsyncCrossingSink_io_out_0_a_bits_data;
  assign dmInner_io_dmi_in_0_d_ready = TLAsyncCrossingSink_io_out_0_d_ready;
  assign dmInner_io_dmactive = _T_164;
  assign dmInner_io_innerCtrl_valid = _T_159_valid;
  assign dmInner_io_innerCtrl_bits_resumereq = _T_159_bits_resumereq;
  assign dmInner_io_innerCtrl_bits_hartsel = _T_159_bits_hartsel;
  assign dmInner_io_debugUnavail_0 = io_debugUnavail_0;
  assign TLAsyncCrossingSink_clock = clock;
  assign TLAsyncCrossingSink_reset = reset;
  assign TLAsyncCrossingSink_io_in_0_a_mem_0_opcode = io_dmi_in_0_a_mem_0_opcode;
  assign TLAsyncCrossingSink_io_in_0_a_mem_0_size = io_dmi_in_0_a_mem_0_size;
  assign TLAsyncCrossingSink_io_in_0_a_mem_0_source = io_dmi_in_0_a_mem_0_source;
  assign TLAsyncCrossingSink_io_in_0_a_mem_0_address = io_dmi_in_0_a_mem_0_address;
  assign TLAsyncCrossingSink_io_in_0_a_mem_0_mask = io_dmi_in_0_a_mem_0_mask;
  assign TLAsyncCrossingSink_io_in_0_a_mem_0_data = io_dmi_in_0_a_mem_0_data;
  assign TLAsyncCrossingSink_io_in_0_a_widx = io_dmi_in_0_a_widx;
  assign TLAsyncCrossingSink_io_in_0_a_widx_valid = io_dmi_in_0_a_widx_valid;
  assign TLAsyncCrossingSink_io_in_0_a_source_reset_n = io_dmi_in_0_a_source_reset_n;
  assign TLAsyncCrossingSink_io_in_0_d_ridx = io_dmi_in_0_d_ridx;
  assign TLAsyncCrossingSink_io_in_0_d_ridx_valid = io_dmi_in_0_d_ridx_valid;
  assign TLAsyncCrossingSink_io_in_0_d_sink_reset_n = io_dmi_in_0_d_sink_reset_n;
  assign TLAsyncCrossingSink_io_out_0_a_ready = dmInner_io_dmi_in_0_a_ready;
  assign TLAsyncCrossingSink_io_out_0_d_valid = dmInner_io_dmi_in_0_d_valid;
  assign TLAsyncCrossingSink_io_out_0_d_bits_opcode = dmInner_io_dmi_in_0_d_bits_opcode;
  assign TLAsyncCrossingSink_io_out_0_d_bits_param = dmInner_io_dmi_in_0_d_bits_param;
  assign TLAsyncCrossingSink_io_out_0_d_bits_size = dmInner_io_dmi_in_0_d_bits_size;
  assign TLAsyncCrossingSink_io_out_0_d_bits_source = dmInner_io_dmi_in_0_d_bits_source;
  assign TLAsyncCrossingSink_io_out_0_d_bits_sink = dmInner_io_dmi_in_0_d_bits_sink;
  assign TLAsyncCrossingSink_io_out_0_d_bits_data = dmInner_io_dmi_in_0_d_bits_data;
  assign TLAsyncCrossingSink_io_out_0_d_bits_error = dmInner_io_dmi_in_0_d_bits_error;
  assign AsyncQueueSink_clock = clock;
  assign AsyncQueueSink_reset = reset;
  assign AsyncQueueSink_io_deq_ready = _T_159_ready;
  assign AsyncQueueSink_io_widx = io_innerCtrl_widx;
  assign AsyncQueueSink_io_mem_0_resumereq = io_innerCtrl_mem_0_resumereq;
  assign AsyncQueueSink_io_mem_0_hartsel = io_innerCtrl_mem_0_hartsel;
  assign AsyncQueueSink_io_source_reset_n = io_innerCtrl_source_reset_n;
  assign AsyncQueueSink_io_widx_valid = io_innerCtrl_widx_valid;
  assign _T_154 = AsyncQueueSink_reset == 1'h0;
  assign _T_159_ready = dmInner_io_innerCtrl_ready;
  assign _T_159_valid = AsyncQueueSink_io_deq_valid;
  assign _T_159_bits_resumereq = AsyncQueueSink_io_deq_bits_resumereq;
  assign _T_159_bits_hartsel = AsyncQueueSink_io_deq_bits_hartsel;
  assign _T_163 = ~ io_dmactive;
  assign ResetCatchAndSync_clock = clock;
  assign ResetCatchAndSync_reset = _T_163;
  assign _T_164 = ~ ResetCatchAndSync_io_sync_reset;
endmodule
module TLDebugModule_debug(
  input         clock,
  input         reset,
  output        io_debugInterrupts_0_0,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [1:0]  io_in_0_a_bits_size,
  input  [9:0]  io_in_0_a_bits_source,
  input  [11:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [1:0]  io_in_0_d_bits_size,
  output [9:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_ctrl_debugUnavail_0,
  output        io_ctrl_ndreset,
  output        io_dmi_dmi_req_ready,
  input         io_dmi_dmi_req_valid,
  input  [6:0]  io_dmi_dmi_req_bits_addr,
  input  [31:0] io_dmi_dmi_req_bits_data,
  input  [1:0]  io_dmi_dmi_req_bits_op,
  input         io_dmi_dmi_resp_ready,
  output        io_dmi_dmi_resp_valid,
  output [31:0] io_dmi_dmi_resp_bits_data,
  output [1:0]  io_dmi_dmi_resp_bits_resp,
  input         io_dmi_dmiClock,
  input         io_dmi_dmiReset
);
  wire  dmOuter_clock;
  wire  dmOuter_reset;
  wire  dmOuter_io_debugInterrupts_0_0;
  wire [2:0] dmOuter_io_dmiInner_0_a_mem_0_opcode;
  wire [1:0] dmOuter_io_dmiInner_0_a_mem_0_size;
  wire  dmOuter_io_dmiInner_0_a_mem_0_source;
  wire [8:0] dmOuter_io_dmiInner_0_a_mem_0_address;
  wire [3:0] dmOuter_io_dmiInner_0_a_mem_0_mask;
  wire [31:0] dmOuter_io_dmiInner_0_a_mem_0_data;
  wire  dmOuter_io_dmiInner_0_a_ridx;
  wire  dmOuter_io_dmiInner_0_a_widx;
  wire  dmOuter_io_dmiInner_0_a_ridx_valid;
  wire  dmOuter_io_dmiInner_0_a_widx_valid;
  wire  dmOuter_io_dmiInner_0_a_source_reset_n;
  wire  dmOuter_io_dmiInner_0_a_sink_reset_n;
  wire [2:0] dmOuter_io_dmiInner_0_d_mem_0_opcode;
  wire [1:0] dmOuter_io_dmiInner_0_d_mem_0_param;
  wire [1:0] dmOuter_io_dmiInner_0_d_mem_0_size;
  wire  dmOuter_io_dmiInner_0_d_mem_0_source;
  wire  dmOuter_io_dmiInner_0_d_mem_0_sink;
  wire [31:0] dmOuter_io_dmiInner_0_d_mem_0_data;
  wire  dmOuter_io_dmiInner_0_d_mem_0_error;
  wire  dmOuter_io_dmiInner_0_d_ridx;
  wire  dmOuter_io_dmiInner_0_d_widx;
  wire  dmOuter_io_dmiInner_0_d_ridx_valid;
  wire  dmOuter_io_dmiInner_0_d_widx_valid;
  wire  dmOuter_io_dmiInner_0_d_source_reset_n;
  wire  dmOuter_io_dmiInner_0_d_sink_reset_n;
  wire  dmOuter_io_dmi_req_ready;
  wire  dmOuter_io_dmi_req_valid;
  wire [6:0] dmOuter_io_dmi_req_bits_addr;
  wire [31:0] dmOuter_io_dmi_req_bits_data;
  wire [1:0] dmOuter_io_dmi_req_bits_op;
  wire  dmOuter_io_dmi_resp_ready;
  wire  dmOuter_io_dmi_resp_valid;
  wire [31:0] dmOuter_io_dmi_resp_bits_data;
  wire [1:0] dmOuter_io_dmi_resp_bits_resp;
  wire  dmOuter_io_ctrl_ndreset;
  wire  dmOuter_io_ctrl_dmactive;
  wire  dmOuter_io_innerCtrl_mem_0_resumereq;
  wire [9:0] dmOuter_io_innerCtrl_mem_0_hartsel;
  wire  dmOuter_io_innerCtrl_ridx;
  wire  dmOuter_io_innerCtrl_widx;
  wire  dmOuter_io_innerCtrl_ridx_valid;
  wire  dmOuter_io_innerCtrl_widx_valid;
  wire  dmOuter_io_innerCtrl_source_reset_n;
  wire  dmOuter_io_innerCtrl_sink_reset_n;
  wire  dmInner_clock;
  wire  dmInner_reset;
  wire [2:0] dmInner_io_dmi_in_0_a_mem_0_opcode;
  wire [1:0] dmInner_io_dmi_in_0_a_mem_0_size;
  wire  dmInner_io_dmi_in_0_a_mem_0_source;
  wire [8:0] dmInner_io_dmi_in_0_a_mem_0_address;
  wire [3:0] dmInner_io_dmi_in_0_a_mem_0_mask;
  wire [31:0] dmInner_io_dmi_in_0_a_mem_0_data;
  wire  dmInner_io_dmi_in_0_a_ridx;
  wire  dmInner_io_dmi_in_0_a_widx;
  wire  dmInner_io_dmi_in_0_a_ridx_valid;
  wire  dmInner_io_dmi_in_0_a_widx_valid;
  wire  dmInner_io_dmi_in_0_a_source_reset_n;
  wire  dmInner_io_dmi_in_0_a_sink_reset_n;
  wire [2:0] dmInner_io_dmi_in_0_d_mem_0_opcode;
  wire [1:0] dmInner_io_dmi_in_0_d_mem_0_param;
  wire [1:0] dmInner_io_dmi_in_0_d_mem_0_size;
  wire  dmInner_io_dmi_in_0_d_mem_0_source;
  wire  dmInner_io_dmi_in_0_d_mem_0_sink;
  wire [31:0] dmInner_io_dmi_in_0_d_mem_0_data;
  wire  dmInner_io_dmi_in_0_d_mem_0_error;
  wire  dmInner_io_dmi_in_0_d_ridx;
  wire  dmInner_io_dmi_in_0_d_widx;
  wire  dmInner_io_dmi_in_0_d_ridx_valid;
  wire  dmInner_io_dmi_in_0_d_widx_valid;
  wire  dmInner_io_dmi_in_0_d_source_reset_n;
  wire  dmInner_io_dmi_in_0_d_sink_reset_n;
  wire  dmInner_io_tl_in_0_a_ready;
  wire  dmInner_io_tl_in_0_a_valid;
  wire [2:0] dmInner_io_tl_in_0_a_bits_opcode;
  wire [1:0] dmInner_io_tl_in_0_a_bits_size;
  wire [9:0] dmInner_io_tl_in_0_a_bits_source;
  wire [11:0] dmInner_io_tl_in_0_a_bits_address;
  wire [3:0] dmInner_io_tl_in_0_a_bits_mask;
  wire [31:0] dmInner_io_tl_in_0_a_bits_data;
  wire  dmInner_io_tl_in_0_d_ready;
  wire  dmInner_io_tl_in_0_d_valid;
  wire [2:0] dmInner_io_tl_in_0_d_bits_opcode;
  wire [1:0] dmInner_io_tl_in_0_d_bits_param;
  wire [1:0] dmInner_io_tl_in_0_d_bits_size;
  wire [9:0] dmInner_io_tl_in_0_d_bits_source;
  wire  dmInner_io_tl_in_0_d_bits_sink;
  wire [31:0] dmInner_io_tl_in_0_d_bits_data;
  wire  dmInner_io_tl_in_0_d_bits_error;
  wire  dmInner_io_dmactive;
  wire  dmInner_io_innerCtrl_mem_0_resumereq;
  wire [9:0] dmInner_io_innerCtrl_mem_0_hartsel;
  wire  dmInner_io_innerCtrl_ridx;
  wire  dmInner_io_innerCtrl_widx;
  wire  dmInner_io_innerCtrl_ridx_valid;
  wire  dmInner_io_innerCtrl_widx_valid;
  wire  dmInner_io_innerCtrl_source_reset_n;
  wire  dmInner_io_innerCtrl_sink_reset_n;
  wire  dmInner_io_debugUnavail_0;
  TLDebugModuleOuterAsync_dmOuter dmOuter (
    .clock(dmOuter_clock),
    .reset(dmOuter_reset),
    .io_debugInterrupts_0_0(dmOuter_io_debugInterrupts_0_0),
    .io_dmiInner_0_a_mem_0_opcode(dmOuter_io_dmiInner_0_a_mem_0_opcode),
    .io_dmiInner_0_a_mem_0_size(dmOuter_io_dmiInner_0_a_mem_0_size),
    .io_dmiInner_0_a_mem_0_source(dmOuter_io_dmiInner_0_a_mem_0_source),
    .io_dmiInner_0_a_mem_0_address(dmOuter_io_dmiInner_0_a_mem_0_address),
    .io_dmiInner_0_a_mem_0_mask(dmOuter_io_dmiInner_0_a_mem_0_mask),
    .io_dmiInner_0_a_mem_0_data(dmOuter_io_dmiInner_0_a_mem_0_data),
    .io_dmiInner_0_a_ridx(dmOuter_io_dmiInner_0_a_ridx),
    .io_dmiInner_0_a_widx(dmOuter_io_dmiInner_0_a_widx),
    .io_dmiInner_0_a_ridx_valid(dmOuter_io_dmiInner_0_a_ridx_valid),
    .io_dmiInner_0_a_widx_valid(dmOuter_io_dmiInner_0_a_widx_valid),
    .io_dmiInner_0_a_source_reset_n(dmOuter_io_dmiInner_0_a_source_reset_n),
    .io_dmiInner_0_a_sink_reset_n(dmOuter_io_dmiInner_0_a_sink_reset_n),
    .io_dmiInner_0_d_mem_0_opcode(dmOuter_io_dmiInner_0_d_mem_0_opcode),
    .io_dmiInner_0_d_mem_0_param(dmOuter_io_dmiInner_0_d_mem_0_param),
    .io_dmiInner_0_d_mem_0_size(dmOuter_io_dmiInner_0_d_mem_0_size),
    .io_dmiInner_0_d_mem_0_source(dmOuter_io_dmiInner_0_d_mem_0_source),
    .io_dmiInner_0_d_mem_0_sink(dmOuter_io_dmiInner_0_d_mem_0_sink),
    .io_dmiInner_0_d_mem_0_data(dmOuter_io_dmiInner_0_d_mem_0_data),
    .io_dmiInner_0_d_mem_0_error(dmOuter_io_dmiInner_0_d_mem_0_error),
    .io_dmiInner_0_d_ridx(dmOuter_io_dmiInner_0_d_ridx),
    .io_dmiInner_0_d_widx(dmOuter_io_dmiInner_0_d_widx),
    .io_dmiInner_0_d_ridx_valid(dmOuter_io_dmiInner_0_d_ridx_valid),
    .io_dmiInner_0_d_widx_valid(dmOuter_io_dmiInner_0_d_widx_valid),
    .io_dmiInner_0_d_source_reset_n(dmOuter_io_dmiInner_0_d_source_reset_n),
    .io_dmiInner_0_d_sink_reset_n(dmOuter_io_dmiInner_0_d_sink_reset_n),
    .io_dmi_req_ready(dmOuter_io_dmi_req_ready),
    .io_dmi_req_valid(dmOuter_io_dmi_req_valid),
    .io_dmi_req_bits_addr(dmOuter_io_dmi_req_bits_addr),
    .io_dmi_req_bits_data(dmOuter_io_dmi_req_bits_data),
    .io_dmi_req_bits_op(dmOuter_io_dmi_req_bits_op),
    .io_dmi_resp_ready(dmOuter_io_dmi_resp_ready),
    .io_dmi_resp_valid(dmOuter_io_dmi_resp_valid),
    .io_dmi_resp_bits_data(dmOuter_io_dmi_resp_bits_data),
    .io_dmi_resp_bits_resp(dmOuter_io_dmi_resp_bits_resp),
    .io_ctrl_ndreset(dmOuter_io_ctrl_ndreset),
    .io_ctrl_dmactive(dmOuter_io_ctrl_dmactive),
    .io_innerCtrl_mem_0_resumereq(dmOuter_io_innerCtrl_mem_0_resumereq),
    .io_innerCtrl_mem_0_hartsel(dmOuter_io_innerCtrl_mem_0_hartsel),
    .io_innerCtrl_ridx(dmOuter_io_innerCtrl_ridx),
    .io_innerCtrl_widx(dmOuter_io_innerCtrl_widx),
    .io_innerCtrl_ridx_valid(dmOuter_io_innerCtrl_ridx_valid),
    .io_innerCtrl_widx_valid(dmOuter_io_innerCtrl_widx_valid),
    .io_innerCtrl_source_reset_n(dmOuter_io_innerCtrl_source_reset_n),
    .io_innerCtrl_sink_reset_n(dmOuter_io_innerCtrl_sink_reset_n)
  );
  TLDebugModuleInnerAsync_dmInner dmInner (
    .clock(dmInner_clock),
    .reset(dmInner_reset),
    .io_dmi_in_0_a_mem_0_opcode(dmInner_io_dmi_in_0_a_mem_0_opcode),
    .io_dmi_in_0_a_mem_0_size(dmInner_io_dmi_in_0_a_mem_0_size),
    .io_dmi_in_0_a_mem_0_source(dmInner_io_dmi_in_0_a_mem_0_source),
    .io_dmi_in_0_a_mem_0_address(dmInner_io_dmi_in_0_a_mem_0_address),
    .io_dmi_in_0_a_mem_0_mask(dmInner_io_dmi_in_0_a_mem_0_mask),
    .io_dmi_in_0_a_mem_0_data(dmInner_io_dmi_in_0_a_mem_0_data),
    .io_dmi_in_0_a_ridx(dmInner_io_dmi_in_0_a_ridx),
    .io_dmi_in_0_a_widx(dmInner_io_dmi_in_0_a_widx),
    .io_dmi_in_0_a_ridx_valid(dmInner_io_dmi_in_0_a_ridx_valid),
    .io_dmi_in_0_a_widx_valid(dmInner_io_dmi_in_0_a_widx_valid),
    .io_dmi_in_0_a_source_reset_n(dmInner_io_dmi_in_0_a_source_reset_n),
    .io_dmi_in_0_a_sink_reset_n(dmInner_io_dmi_in_0_a_sink_reset_n),
    .io_dmi_in_0_d_mem_0_opcode(dmInner_io_dmi_in_0_d_mem_0_opcode),
    .io_dmi_in_0_d_mem_0_param(dmInner_io_dmi_in_0_d_mem_0_param),
    .io_dmi_in_0_d_mem_0_size(dmInner_io_dmi_in_0_d_mem_0_size),
    .io_dmi_in_0_d_mem_0_source(dmInner_io_dmi_in_0_d_mem_0_source),
    .io_dmi_in_0_d_mem_0_sink(dmInner_io_dmi_in_0_d_mem_0_sink),
    .io_dmi_in_0_d_mem_0_data(dmInner_io_dmi_in_0_d_mem_0_data),
    .io_dmi_in_0_d_mem_0_error(dmInner_io_dmi_in_0_d_mem_0_error),
    .io_dmi_in_0_d_ridx(dmInner_io_dmi_in_0_d_ridx),
    .io_dmi_in_0_d_widx(dmInner_io_dmi_in_0_d_widx),
    .io_dmi_in_0_d_ridx_valid(dmInner_io_dmi_in_0_d_ridx_valid),
    .io_dmi_in_0_d_widx_valid(dmInner_io_dmi_in_0_d_widx_valid),
    .io_dmi_in_0_d_source_reset_n(dmInner_io_dmi_in_0_d_source_reset_n),
    .io_dmi_in_0_d_sink_reset_n(dmInner_io_dmi_in_0_d_sink_reset_n),
    .io_tl_in_0_a_ready(dmInner_io_tl_in_0_a_ready),
    .io_tl_in_0_a_valid(dmInner_io_tl_in_0_a_valid),
    .io_tl_in_0_a_bits_opcode(dmInner_io_tl_in_0_a_bits_opcode),
    .io_tl_in_0_a_bits_size(dmInner_io_tl_in_0_a_bits_size),
    .io_tl_in_0_a_bits_source(dmInner_io_tl_in_0_a_bits_source),
    .io_tl_in_0_a_bits_address(dmInner_io_tl_in_0_a_bits_address),
    .io_tl_in_0_a_bits_mask(dmInner_io_tl_in_0_a_bits_mask),
    .io_tl_in_0_a_bits_data(dmInner_io_tl_in_0_a_bits_data),
    .io_tl_in_0_d_ready(dmInner_io_tl_in_0_d_ready),
    .io_tl_in_0_d_valid(dmInner_io_tl_in_0_d_valid),
    .io_tl_in_0_d_bits_opcode(dmInner_io_tl_in_0_d_bits_opcode),
    .io_tl_in_0_d_bits_param(dmInner_io_tl_in_0_d_bits_param),
    .io_tl_in_0_d_bits_size(dmInner_io_tl_in_0_d_bits_size),
    .io_tl_in_0_d_bits_source(dmInner_io_tl_in_0_d_bits_source),
    .io_tl_in_0_d_bits_sink(dmInner_io_tl_in_0_d_bits_sink),
    .io_tl_in_0_d_bits_data(dmInner_io_tl_in_0_d_bits_data),
    .io_tl_in_0_d_bits_error(dmInner_io_tl_in_0_d_bits_error),
    .io_dmactive(dmInner_io_dmactive),
    .io_innerCtrl_mem_0_resumereq(dmInner_io_innerCtrl_mem_0_resumereq),
    .io_innerCtrl_mem_0_hartsel(dmInner_io_innerCtrl_mem_0_hartsel),
    .io_innerCtrl_ridx(dmInner_io_innerCtrl_ridx),
    .io_innerCtrl_widx(dmInner_io_innerCtrl_widx),
    .io_innerCtrl_ridx_valid(dmInner_io_innerCtrl_ridx_valid),
    .io_innerCtrl_widx_valid(dmInner_io_innerCtrl_widx_valid),
    .io_innerCtrl_source_reset_n(dmInner_io_innerCtrl_source_reset_n),
    .io_innerCtrl_sink_reset_n(dmInner_io_innerCtrl_sink_reset_n),
    .io_debugUnavail_0(dmInner_io_debugUnavail_0)
  );
  assign io_debugInterrupts_0_0 = dmOuter_io_debugInterrupts_0_0;
  assign io_in_0_a_ready = dmInner_io_tl_in_0_a_ready;
  assign io_in_0_d_valid = dmInner_io_tl_in_0_d_valid;
  assign io_in_0_d_bits_opcode = dmInner_io_tl_in_0_d_bits_opcode;
  assign io_in_0_d_bits_param = dmInner_io_tl_in_0_d_bits_param;
  assign io_in_0_d_bits_size = dmInner_io_tl_in_0_d_bits_size;
  assign io_in_0_d_bits_source = dmInner_io_tl_in_0_d_bits_source;
  assign io_in_0_d_bits_sink = dmInner_io_tl_in_0_d_bits_sink;
  assign io_in_0_d_bits_data = dmInner_io_tl_in_0_d_bits_data;
  assign io_in_0_d_bits_error = dmInner_io_tl_in_0_d_bits_error;
  assign io_ctrl_ndreset = dmOuter_io_ctrl_ndreset;
  assign io_dmi_dmi_req_ready = dmOuter_io_dmi_req_ready;
  assign io_dmi_dmi_resp_valid = dmOuter_io_dmi_resp_valid;
  assign io_dmi_dmi_resp_bits_data = dmOuter_io_dmi_resp_bits_data;
  assign io_dmi_dmi_resp_bits_resp = dmOuter_io_dmi_resp_bits_resp;
  assign dmOuter_clock = io_dmi_dmiClock;
  assign dmOuter_reset = io_dmi_dmiReset;
  assign dmOuter_io_dmiInner_0_a_ridx = dmInner_io_dmi_in_0_a_ridx;
  assign dmOuter_io_dmiInner_0_a_ridx_valid = dmInner_io_dmi_in_0_a_ridx_valid;
  assign dmOuter_io_dmiInner_0_a_sink_reset_n = dmInner_io_dmi_in_0_a_sink_reset_n;
  assign dmOuter_io_dmiInner_0_d_mem_0_opcode = dmInner_io_dmi_in_0_d_mem_0_opcode;
  assign dmOuter_io_dmiInner_0_d_mem_0_param = dmInner_io_dmi_in_0_d_mem_0_param;
  assign dmOuter_io_dmiInner_0_d_mem_0_size = dmInner_io_dmi_in_0_d_mem_0_size;
  assign dmOuter_io_dmiInner_0_d_mem_0_source = dmInner_io_dmi_in_0_d_mem_0_source;
  assign dmOuter_io_dmiInner_0_d_mem_0_sink = dmInner_io_dmi_in_0_d_mem_0_sink;
  assign dmOuter_io_dmiInner_0_d_mem_0_data = dmInner_io_dmi_in_0_d_mem_0_data;
  assign dmOuter_io_dmiInner_0_d_mem_0_error = dmInner_io_dmi_in_0_d_mem_0_error;
  assign dmOuter_io_dmiInner_0_d_widx = dmInner_io_dmi_in_0_d_widx;
  assign dmOuter_io_dmiInner_0_d_widx_valid = dmInner_io_dmi_in_0_d_widx_valid;
  assign dmOuter_io_dmiInner_0_d_source_reset_n = dmInner_io_dmi_in_0_d_source_reset_n;
  assign dmOuter_io_dmi_req_valid = io_dmi_dmi_req_valid;
  assign dmOuter_io_dmi_req_bits_addr = io_dmi_dmi_req_bits_addr;
  assign dmOuter_io_dmi_req_bits_data = io_dmi_dmi_req_bits_data;
  assign dmOuter_io_dmi_req_bits_op = io_dmi_dmi_req_bits_op;
  assign dmOuter_io_dmi_resp_ready = io_dmi_dmi_resp_ready;
  assign dmOuter_io_innerCtrl_ridx = dmInner_io_innerCtrl_ridx;
  assign dmOuter_io_innerCtrl_ridx_valid = dmInner_io_innerCtrl_ridx_valid;
  assign dmOuter_io_innerCtrl_sink_reset_n = dmInner_io_innerCtrl_sink_reset_n;
  assign dmInner_clock = clock;
  assign dmInner_reset = reset;
  assign dmInner_io_dmi_in_0_a_mem_0_opcode = dmOuter_io_dmiInner_0_a_mem_0_opcode;
  assign dmInner_io_dmi_in_0_a_mem_0_size = dmOuter_io_dmiInner_0_a_mem_0_size;
  assign dmInner_io_dmi_in_0_a_mem_0_source = dmOuter_io_dmiInner_0_a_mem_0_source;
  assign dmInner_io_dmi_in_0_a_mem_0_address = dmOuter_io_dmiInner_0_a_mem_0_address;
  assign dmInner_io_dmi_in_0_a_mem_0_mask = dmOuter_io_dmiInner_0_a_mem_0_mask;
  assign dmInner_io_dmi_in_0_a_mem_0_data = dmOuter_io_dmiInner_0_a_mem_0_data;
  assign dmInner_io_dmi_in_0_a_widx = dmOuter_io_dmiInner_0_a_widx;
  assign dmInner_io_dmi_in_0_a_widx_valid = dmOuter_io_dmiInner_0_a_widx_valid;
  assign dmInner_io_dmi_in_0_a_source_reset_n = dmOuter_io_dmiInner_0_a_source_reset_n;
  assign dmInner_io_dmi_in_0_d_ridx = dmOuter_io_dmiInner_0_d_ridx;
  assign dmInner_io_dmi_in_0_d_ridx_valid = dmOuter_io_dmiInner_0_d_ridx_valid;
  assign dmInner_io_dmi_in_0_d_sink_reset_n = dmOuter_io_dmiInner_0_d_sink_reset_n;
  assign dmInner_io_tl_in_0_a_valid = io_in_0_a_valid;
  assign dmInner_io_tl_in_0_a_bits_opcode = io_in_0_a_bits_opcode;
  assign dmInner_io_tl_in_0_a_bits_size = io_in_0_a_bits_size;
  assign dmInner_io_tl_in_0_a_bits_source = io_in_0_a_bits_source;
  assign dmInner_io_tl_in_0_a_bits_address = io_in_0_a_bits_address;
  assign dmInner_io_tl_in_0_a_bits_mask = io_in_0_a_bits_mask;
  assign dmInner_io_tl_in_0_a_bits_data = io_in_0_a_bits_data;
  assign dmInner_io_tl_in_0_d_ready = io_in_0_d_ready;
  assign dmInner_io_dmactive = dmOuter_io_ctrl_dmactive;
  assign dmInner_io_innerCtrl_mem_0_resumereq = dmOuter_io_innerCtrl_mem_0_resumereq;
  assign dmInner_io_innerCtrl_mem_0_hartsel = dmOuter_io_innerCtrl_mem_0_hartsel;
  assign dmInner_io_innerCtrl_widx = dmOuter_io_innerCtrl_widx;
  assign dmInner_io_innerCtrl_widx_valid = dmOuter_io_innerCtrl_widx_valid;
  assign dmInner_io_innerCtrl_source_reset_n = dmOuter_io_innerCtrl_source_reset_n;
  assign dmInner_io_debugUnavail_0 = io_ctrl_debugUnavail_0;
endmodule
module TLXbar_tileBus(
  input         clock,
  input         reset,
  output        io_in_1_a_ready,
  input         io_in_1_a_valid,
  input  [2:0]  io_in_1_a_bits_opcode,
  input  [2:0]  io_in_1_a_bits_param,
  input  [3:0]  io_in_1_a_bits_size,
  input         io_in_1_a_bits_source,
  input  [31:0] io_in_1_a_bits_address,
  input  [3:0]  io_in_1_a_bits_mask,
  input  [31:0] io_in_1_a_bits_data,
  input         io_in_1_d_ready,
  output        io_in_1_d_valid,
  output [2:0]  io_in_1_d_bits_opcode,
  output [3:0]  io_in_1_d_bits_size,
  output [31:0] io_in_1_d_bits_data,
  output        io_in_1_d_bits_error,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  output        io_in_0_b_valid,
  output [1:0]  io_in_0_b_bits_param,
  output [31:0] io_in_0_b_bits_address,
  output        io_in_0_c_ready,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output        io_in_0_d_bits_source,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_e_ready,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input         io_out_0_d_bits_source,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  _T_900;
  wire [26:0] _T_1036;
  wire [11:0] _T_1037;
  wire [11:0] _T_1038;
  wire [9:0] _T_1039;
  wire  _T_1040;
  wire  _T_1042;
  wire [9:0] _T_1044;
  wire [26:0] _T_1047;
  wire [11:0] _T_1048;
  wire [11:0] _T_1049;
  wire [9:0] _T_1050;
  wire  _T_1051;
  wire  _T_1053;
  wire [9:0] _T_1055;
  wire  _T_1305;
  wire  _T_1306;
  wire  _T_1309;
  wire  _T_1311;
  wire  _T_1312;
  reg [9:0] _T_1367;
  reg [31:0] _RAND_0;
  wire  _T_1369;
  wire  _T_1370;
  wire [1:0] _T_1371;
  wire  _T_1373;
  wire  _T_1374;
  wire  _T_1376;
  reg [1:0] _T_1380;
  reg [31:0] _RAND_1;
  wire [1:0] _T_1381;
  wire [1:0] _T_1382;
  wire [3:0] _T_1383;
  wire [2:0] _T_1384;
  wire [3:0] _GEN_1;
  wire [3:0] _T_1385;
  wire [2:0] _T_1387;
  wire [3:0] _GEN_2;
  wire [3:0] _T_1388;
  wire [3:0] _GEN_3;
  wire [3:0] _T_1389;
  wire [1:0] _T_1390;
  wire [1:0] _T_1391;
  wire [1:0] _T_1392;
  wire [1:0] _T_1393;
  wire  _T_1395;
  wire  _T_1396;
  wire [1:0] _T_1397;
  wire [2:0] _GEN_4;
  wire [2:0] _T_1398;
  wire [1:0] _T_1399;
  wire [1:0] _T_1400;
  wire [1:0] _GEN_0;
  wire  _T_1403;
  wire  _T_1404;
  wire  _T_1412;
  wire  _T_1413;
  wire  _T_1423;
  wire  _T_1427;
  wire  _T_1432;
  wire  _T_1433;
  wire  _T_1435;
  wire  _T_1437;
  wire  _T_1438;
  wire  _T_1440;
  wire  _T_1442;
  wire  _T_1443;
  wire  _T_1445;
  wire [9:0] _T_1447;
  wire [9:0] _T_1449;
  wire [9:0] _T_1450;
  wire  _T_1451;
  wire [9:0] _GEN_5;
  wire [10:0] _T_1452;
  wire [10:0] _T_1453;
  wire [9:0] _T_1454;
  wire [9:0] _T_1455;
  reg  _T_1473_0;
  reg [31:0] _RAND_2;
  reg  _T_1473_1;
  reg [31:0] _RAND_3;
  wire  _T_1484_0;
  wire  _T_1484_1;
  wire  _T_1492_0;
  wire  _T_1492_1;
  wire  _T_1500;
  wire  _T_1501;
  wire  _T_1505;
  wire  _T_1507;
  wire  _T_1508;
  wire  _T_1511;
  wire [35:0] _T_1513;
  wire [67:0] _T_1514;
  wire [4:0] _T_1515;
  wire [5:0] _T_1516;
  wire [10:0] _T_1517;
  wire [78:0] _T_1518;
  wire [78:0] _T_1520;
  wire [35:0] _T_1521;
  wire [67:0] _T_1522;
  wire [4:0] _T_1523;
  wire [5:0] _T_1524;
  wire [10:0] _T_1525;
  wire [78:0] _T_1526;
  wire [78:0] _T_1528;
  wire [78:0] _T_1529;
  wire [31:0] _T_1534;
  wire [3:0] _T_1535;
  wire [31:0] _T_1536;
  wire  _T_1537;
  wire [3:0] _T_1538;
  wire [2:0] _T_1539;
  wire [2:0] _T_1540;
  wire  _T_1570;
  wire  _T_1577;
  wire  _T_1578;
  wire  _T_1580;
  wire  _T_1643;
  wire  _T_1650;
  wire  _T_1651;
  wire  _T_1653;
  assign io_in_1_a_ready = _T_1501;
  assign io_in_1_d_valid = _T_1306;
  assign io_in_1_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_1_d_bits_size = io_out_0_d_bits_size;
  assign io_in_1_d_bits_data = io_out_0_d_bits_data;
  assign io_in_1_d_bits_error = io_out_0_d_bits_error;
  assign io_in_0_a_ready = _T_1500;
  assign io_in_0_b_valid = 1'h0;
  assign io_in_0_b_bits_param = 2'h0;
  assign io_in_0_b_bits_address = 32'h0;
  assign io_in_0_c_ready = 1'h1;
  assign io_in_0_d_valid = _T_1305;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = 1'h0;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_e_ready = 1'h1;
  assign io_out_0_a_valid = _T_1511;
  assign io_out_0_a_bits_opcode = _T_1540;
  assign io_out_0_a_bits_param = _T_1539;
  assign io_out_0_a_bits_size = _T_1538;
  assign io_out_0_a_bits_source = _T_1537;
  assign io_out_0_a_bits_address = _T_1536;
  assign io_out_0_a_bits_mask = _T_1535;
  assign io_out_0_a_bits_data = _T_1534;
  assign io_out_0_d_ready = _T_1312;
  assign _T_900 = io_out_0_d_bits_source == 1'h0;
  assign _T_1036 = 27'hfff << io_in_0_a_bits_size;
  assign _T_1037 = _T_1036[11:0];
  assign _T_1038 = ~ _T_1037;
  assign _T_1039 = _T_1038[11:2];
  assign _T_1040 = io_in_0_a_bits_opcode[2];
  assign _T_1042 = _T_1040 == 1'h0;
  assign _T_1044 = _T_1042 ? _T_1039 : 10'h0;
  assign _T_1047 = 27'hfff << io_in_1_a_bits_size;
  assign _T_1048 = _T_1047[11:0];
  assign _T_1049 = ~ _T_1048;
  assign _T_1050 = _T_1049[11:2];
  assign _T_1051 = io_in_1_a_bits_opcode[2];
  assign _T_1053 = _T_1051 == 1'h0;
  assign _T_1055 = _T_1053 ? _T_1050 : 10'h0;
  assign _T_1305 = io_out_0_d_valid & io_out_0_d_bits_source;
  assign _T_1306 = io_out_0_d_valid & _T_900;
  assign _T_1309 = io_out_0_d_bits_source ? io_in_0_d_ready : 1'h0;
  assign _T_1311 = _T_900 ? io_in_1_d_ready : 1'h0;
  assign _T_1312 = _T_1309 | _T_1311;
  assign _T_1369 = _T_1367 == 10'h0;
  assign _T_1370 = _T_1369 & io_out_0_a_ready;
  assign _T_1371 = {io_in_1_a_valid,io_in_0_a_valid};
  assign _T_1373 = _T_1371 == _T_1371;
  assign _T_1374 = _T_1373 | reset;
  assign _T_1376 = _T_1374 == 1'h0;
  assign _T_1381 = ~ _T_1380;
  assign _T_1382 = _T_1371 & _T_1381;
  assign _T_1383 = {_T_1382,_T_1371};
  assign _T_1384 = _T_1383[3:1];
  assign _GEN_1 = {{1'd0}, _T_1384};
  assign _T_1385 = _T_1383 | _GEN_1;
  assign _T_1387 = _T_1385[3:1];
  assign _GEN_2 = {{2'd0}, _T_1380};
  assign _T_1388 = _GEN_2 << 2;
  assign _GEN_3 = {{1'd0}, _T_1387};
  assign _T_1389 = _GEN_3 | _T_1388;
  assign _T_1390 = _T_1389[3:2];
  assign _T_1391 = _T_1389[1:0];
  assign _T_1392 = _T_1390 & _T_1391;
  assign _T_1393 = ~ _T_1392;
  assign _T_1395 = _T_1371 != 2'h0;
  assign _T_1396 = _T_1370 & _T_1395;
  assign _T_1397 = _T_1393 & _T_1371;
  assign _GEN_4 = {{1'd0}, _T_1397};
  assign _T_1398 = _GEN_4 << 1;
  assign _T_1399 = _T_1398[1:0];
  assign _T_1400 = _T_1397 | _T_1399;
  assign _GEN_0 = _T_1396 ? _T_1400 : _T_1380;
  assign _T_1403 = _T_1393[0];
  assign _T_1404 = _T_1393[1];
  assign _T_1412 = _T_1403 & io_in_0_a_valid;
  assign _T_1413 = _T_1404 & io_in_1_a_valid;
  assign _T_1423 = _T_1412 | _T_1413;
  assign _T_1427 = _T_1412 == 1'h0;
  assign _T_1432 = _T_1413 == 1'h0;
  assign _T_1433 = _T_1427 | _T_1432;
  assign _T_1435 = _T_1433 | reset;
  assign _T_1437 = _T_1435 == 1'h0;
  assign _T_1438 = io_in_0_a_valid | io_in_1_a_valid;
  assign _T_1440 = _T_1438 == 1'h0;
  assign _T_1442 = _T_1440 | _T_1423;
  assign _T_1443 = _T_1442 | reset;
  assign _T_1445 = _T_1443 == 1'h0;
  assign _T_1447 = _T_1412 ? _T_1044 : 10'h0;
  assign _T_1449 = _T_1413 ? _T_1055 : 10'h0;
  assign _T_1450 = _T_1447 | _T_1449;
  assign _T_1451 = io_out_0_a_ready & _T_1511;
  assign _GEN_5 = {{9'd0}, _T_1451};
  assign _T_1452 = _T_1367 - _GEN_5;
  assign _T_1453 = $unsigned(_T_1452);
  assign _T_1454 = _T_1453[9:0];
  assign _T_1455 = _T_1370 ? _T_1450 : _T_1454;
  assign _T_1484_0 = _T_1369 ? _T_1412 : _T_1473_0;
  assign _T_1484_1 = _T_1369 ? _T_1413 : _T_1473_1;
  assign _T_1492_0 = _T_1369 ? _T_1403 : _T_1473_0;
  assign _T_1492_1 = _T_1369 ? _T_1404 : _T_1473_1;
  assign _T_1500 = io_out_0_a_ready & _T_1492_0;
  assign _T_1501 = io_out_0_a_ready & _T_1492_1;
  assign _T_1505 = _T_1473_0 ? io_in_0_a_valid : 1'h0;
  assign _T_1507 = _T_1473_1 ? io_in_1_a_valid : 1'h0;
  assign _T_1508 = _T_1505 | _T_1507;
  assign _T_1511 = _T_1369 ? _T_1438 : _T_1508;
  assign _T_1513 = {io_in_0_a_bits_address,io_in_0_a_bits_mask};
  assign _T_1514 = {_T_1513,io_in_0_a_bits_data};
  assign _T_1515 = {io_in_0_a_bits_size,1'h1};
  assign _T_1516 = {io_in_0_a_bits_opcode,io_in_0_a_bits_param};
  assign _T_1517 = {_T_1516,_T_1515};
  assign _T_1518 = {_T_1517,_T_1514};
  assign _T_1520 = _T_1484_0 ? _T_1518 : 79'h0;
  assign _T_1521 = {io_in_1_a_bits_address,io_in_1_a_bits_mask};
  assign _T_1522 = {_T_1521,io_in_1_a_bits_data};
  assign _T_1523 = {io_in_1_a_bits_size,io_in_1_a_bits_source};
  assign _T_1524 = {io_in_1_a_bits_opcode,io_in_1_a_bits_param};
  assign _T_1525 = {_T_1524,_T_1523};
  assign _T_1526 = {_T_1525,_T_1522};
  assign _T_1528 = _T_1484_1 ? _T_1526 : 79'h0;
  assign _T_1529 = _T_1520 | _T_1528;
  assign _T_1534 = _T_1529[31:0];
  assign _T_1535 = _T_1529[35:32];
  assign _T_1536 = _T_1529[67:36];
  assign _T_1537 = _T_1529[68];
  assign _T_1538 = _T_1529[72:69];
  assign _T_1539 = _T_1529[75:73];
  assign _T_1540 = _T_1529[78:76];
  assign _T_1570 = _T_1305 == 1'h0;
  assign _T_1577 = _T_1570 | _T_1305;
  assign _T_1578 = _T_1577 | reset;
  assign _T_1580 = _T_1578 == 1'h0;
  assign _T_1643 = _T_1306 == 1'h0;
  assign _T_1650 = _T_1643 | _T_1306;
  assign _T_1651 = _T_1650 | reset;
  assign _T_1653 = _T_1651 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_1367 = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_1380 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_1473_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_1473_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1367 <= 10'h0;
    end else begin
      if (_T_1370) begin
        _T_1367 <= _T_1450;
      end else begin
        _T_1367 <= _T_1454;
      end
    end
    if (reset) begin
      _T_1380 <= 2'h3;
    end else begin
      if (_T_1396) begin
        _T_1380 <= _T_1400;
      end
    end
    if (reset) begin
      _T_1473_0 <= 1'h0;
    end else begin
      if (_T_1369) begin
        _T_1473_0 <= _T_1412;
      end
    end
    if (reset) begin
      _T_1473_1 <= 1'h0;
    end else begin
      if (_T_1369) begin
        _T_1473_1 <= _T_1413;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1376) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1376) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1437) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1437) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1445) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1445) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1580) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1580) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1653) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1653) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter(
  input        io_in_0_valid,
  input        io_in_0_bits_write,
  input  [7:0] io_in_0_bits_idx,
  input        io_in_1_valid,
  input        io_in_1_bits_write,
  input  [7:0] io_in_1_bits_idx,
  input        io_in_2_valid,
  input        io_in_2_bits_write,
  input  [7:0] io_in_2_bits_idx,
  output       io_in_3_ready,
  input        io_in_3_valid,
  input        io_in_3_bits_write,
  input  [7:0] io_in_3_bits_idx,
  output       io_in_4_ready,
  input        io_in_4_valid,
  input        io_in_4_bits_write,
  input  [7:0] io_in_4_bits_idx,
  output       io_in_5_ready,
  input        io_in_5_valid,
  input        io_in_5_bits_write,
  input  [7:0] io_in_5_bits_idx,
  output       io_in_6_ready,
  input        io_in_6_valid,
  input        io_in_6_bits_write,
  input  [7:0] io_in_6_bits_idx,
  output       io_in_7_ready,
  input        io_in_7_valid,
  input        io_in_7_bits_write,
  input  [7:0] io_in_7_bits_idx,
  input        io_out_ready,
  output       io_out_valid,
  output       io_out_bits_write,
  output [7:0] io_out_bits_idx
);
  wire  _GEN_1;
  wire [7:0] _GEN_2;
  wire  _GEN_7;
  wire [7:0] _GEN_8;
  wire  _GEN_13;
  wire [7:0] _GEN_14;
  wire  _GEN_19;
  wire [7:0] _GEN_20;
  wire  _GEN_25;
  wire [7:0] _GEN_26;
  wire  _GEN_31;
  wire [7:0] _GEN_32;
  wire  _GEN_37;
  wire [7:0] _GEN_38;
  wire  _T_112;
  wire  _T_113;
  wire  _T_114;
  wire  _T_115;
  wire  _T_116;
  wire  _T_117;
  wire  _T_123;
  wire  _T_125;
  wire  _T_127;
  wire  _T_129;
  wire  _T_131;
  wire  _T_135;
  wire  _T_136;
  wire  _T_137;
  wire  _T_138;
  wire  _T_139;
  wire  _T_141;
  wire  _T_142;
  assign io_in_3_ready = _T_135;
  assign io_in_4_ready = _T_136;
  assign io_in_5_ready = _T_137;
  assign io_in_6_ready = _T_138;
  assign io_in_7_ready = _T_139;
  assign io_out_valid = _T_142;
  assign io_out_bits_write = _GEN_37;
  assign io_out_bits_idx = _GEN_38;
  assign _GEN_1 = io_in_6_valid ? io_in_6_bits_write : io_in_7_bits_write;
  assign _GEN_2 = io_in_6_valid ? io_in_6_bits_idx : io_in_7_bits_idx;
  assign _GEN_7 = io_in_5_valid ? io_in_5_bits_write : _GEN_1;
  assign _GEN_8 = io_in_5_valid ? io_in_5_bits_idx : _GEN_2;
  assign _GEN_13 = io_in_4_valid ? io_in_4_bits_write : _GEN_7;
  assign _GEN_14 = io_in_4_valid ? io_in_4_bits_idx : _GEN_8;
  assign _GEN_19 = io_in_3_valid ? io_in_3_bits_write : _GEN_13;
  assign _GEN_20 = io_in_3_valid ? io_in_3_bits_idx : _GEN_14;
  assign _GEN_25 = io_in_2_valid ? io_in_2_bits_write : _GEN_19;
  assign _GEN_26 = io_in_2_valid ? io_in_2_bits_idx : _GEN_20;
  assign _GEN_31 = io_in_1_valid ? io_in_1_bits_write : _GEN_25;
  assign _GEN_32 = io_in_1_valid ? io_in_1_bits_idx : _GEN_26;
  assign _GEN_37 = io_in_0_valid ? io_in_0_bits_write : _GEN_31;
  assign _GEN_38 = io_in_0_valid ? io_in_0_bits_idx : _GEN_32;
  assign _T_112 = io_in_0_valid | io_in_1_valid;
  assign _T_113 = _T_112 | io_in_2_valid;
  assign _T_114 = _T_113 | io_in_3_valid;
  assign _T_115 = _T_114 | io_in_4_valid;
  assign _T_116 = _T_115 | io_in_5_valid;
  assign _T_117 = _T_116 | io_in_6_valid;
  assign _T_123 = _T_113 == 1'h0;
  assign _T_125 = _T_114 == 1'h0;
  assign _T_127 = _T_115 == 1'h0;
  assign _T_129 = _T_116 == 1'h0;
  assign _T_131 = _T_117 == 1'h0;
  assign _T_135 = _T_123 & io_out_ready;
  assign _T_136 = _T_125 & io_out_ready;
  assign _T_137 = _T_127 & io_out_ready;
  assign _T_138 = _T_129 & io_out_ready;
  assign _T_139 = _T_131 & io_out_ready;
  assign _T_141 = _T_131 == 1'h0;
  assign _T_142 = _T_141 | io_in_7_valid;
endmodule
module DCacheDataArray(
  input         clock,
  input         io_req_valid,
  input  [13:0] io_req_bits_addr,
  input         io_req_bits_write,
  input  [31:0] io_req_bits_wdata,
  input  [3:0]  io_req_bits_eccMask,
  output [31:0] io_resp_0
);
  wire  eccMask_0;
  wire  eccMask_1;
  wire  eccMask_2;
  wire  eccMask_3;
  wire [11:0] addr;
  wire [11:0] data_arrays_0_RW0_addr;
  wire  data_arrays_0_RW0_en;
  wire  data_arrays_0_RW0_clk;
  wire  data_arrays_0_RW0_wmode;
  wire [7:0] data_arrays_0_RW0_wdata_0;
  wire [7:0] data_arrays_0_RW0_wdata_1;
  wire [7:0] data_arrays_0_RW0_wdata_2;
  wire [7:0] data_arrays_0_RW0_wdata_3;
  wire [7:0] data_arrays_0_RW0_rdata_0;
  wire [7:0] data_arrays_0_RW0_rdata_1;
  wire [7:0] data_arrays_0_RW0_rdata_2;
  wire [7:0] data_arrays_0_RW0_rdata_3;
  wire  data_arrays_0_RW0_wmask_0;
  wire  data_arrays_0_RW0_wmask_1;
  wire  data_arrays_0_RW0_wmask_2;
  wire  data_arrays_0_RW0_wmask_3;
  wire  _T_28;
  wire [7:0] _T_29;
  wire [7:0] _T_30;
  wire [7:0] _T_31;
  wire [7:0] _T_32;
  wire  _GEN_12;
  wire  _GEN_14;
  wire  _GEN_16;
  wire  _GEN_18;
  wire  _T_55;
  wire  _T_56;
  wire [15:0] _T_74;
  wire [15:0] _T_75;
  wire [31:0] rdata_0_0;
  data_arrays_0 data_arrays_0 (
    .RW0_addr(data_arrays_0_RW0_addr),
    .RW0_en(data_arrays_0_RW0_en),
    .RW0_clk(data_arrays_0_RW0_clk),
    .RW0_wmode(data_arrays_0_RW0_wmode),
    .RW0_wdata_0(data_arrays_0_RW0_wdata_0),
    .RW0_wdata_1(data_arrays_0_RW0_wdata_1),
    .RW0_wdata_2(data_arrays_0_RW0_wdata_2),
    .RW0_wdata_3(data_arrays_0_RW0_wdata_3),
    .RW0_rdata_0(data_arrays_0_RW0_rdata_0),
    .RW0_rdata_1(data_arrays_0_RW0_rdata_1),
    .RW0_rdata_2(data_arrays_0_RW0_rdata_2),
    .RW0_rdata_3(data_arrays_0_RW0_rdata_3),
    .RW0_wmask_0(data_arrays_0_RW0_wmask_0),
    .RW0_wmask_1(data_arrays_0_RW0_wmask_1),
    .RW0_wmask_2(data_arrays_0_RW0_wmask_2),
    .RW0_wmask_3(data_arrays_0_RW0_wmask_3)
  );
  assign io_resp_0 = rdata_0_0;
  assign eccMask_0 = io_req_bits_eccMask[0];
  assign eccMask_1 = io_req_bits_eccMask[1];
  assign eccMask_2 = io_req_bits_eccMask[2];
  assign eccMask_3 = io_req_bits_eccMask[3];
  assign addr = io_req_bits_addr[13:2];
  assign data_arrays_0_RW0_addr = addr;
  assign data_arrays_0_RW0_en = _T_56 | _T_28;
  assign data_arrays_0_RW0_clk = clock;
  assign data_arrays_0_RW0_wmode = _T_28;
  assign data_arrays_0_RW0_wdata_0 = _T_29;
  assign data_arrays_0_RW0_wdata_1 = _T_30;
  assign data_arrays_0_RW0_wdata_2 = _T_31;
  assign data_arrays_0_RW0_wdata_3 = _T_32;
  assign data_arrays_0_RW0_wmask_0 = _GEN_12;
  assign data_arrays_0_RW0_wmask_1 = _GEN_14;
  assign data_arrays_0_RW0_wmask_2 = _GEN_16;
  assign data_arrays_0_RW0_wmask_3 = _GEN_18;
  assign _T_28 = io_req_valid & io_req_bits_write;
  assign _T_29 = io_req_bits_wdata[7:0];
  assign _T_30 = io_req_bits_wdata[15:8];
  assign _T_31 = io_req_bits_wdata[23:16];
  assign _T_32 = io_req_bits_wdata[31:24];
  assign _GEN_12 = _T_28 ? eccMask_0 : 1'h0;
  assign _GEN_14 = _T_28 ? eccMask_1 : 1'h0;
  assign _GEN_16 = _T_28 ? eccMask_2 : 1'h0;
  assign _GEN_18 = _T_28 ? eccMask_3 : 1'h0;
  assign _T_55 = io_req_bits_write == 1'h0;
  assign _T_56 = io_req_valid & _T_55;
  assign _T_74 = {data_arrays_0_RW0_rdata_1,data_arrays_0_RW0_rdata_0};
  assign _T_75 = {data_arrays_0_RW0_rdata_3,data_arrays_0_RW0_rdata_2};
  assign rdata_0_0 = {_T_75,_T_74};
endmodule
module Arbiter_1(
  input         io_in_0_valid,
  input  [13:0] io_in_0_bits_addr,
  input         io_in_0_bits_write,
  input  [31:0] io_in_0_bits_wdata,
  input  [3:0]  io_in_0_bits_eccMask,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [13:0] io_in_1_bits_addr,
  input         io_in_1_bits_write,
  input  [31:0] io_in_1_bits_wdata,
  input  [3:0]  io_in_1_bits_eccMask,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [13:0] io_in_2_bits_addr,
  input         io_in_2_bits_write,
  input  [31:0] io_in_2_bits_wdata,
  input  [3:0]  io_in_2_bits_eccMask,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [13:0] io_in_3_bits_addr,
  input         io_in_3_bits_write,
  input  [31:0] io_in_3_bits_wdata,
  input  [3:0]  io_in_3_bits_eccMask,
  input         io_out_ready,
  output        io_out_valid,
  output [13:0] io_out_bits_addr,
  output        io_out_bits_write,
  output [31:0] io_out_bits_wdata,
  output [3:0]  io_out_bits_eccMask
);
  wire [13:0] _GEN_1;
  wire  _GEN_2;
  wire [31:0] _GEN_3;
  wire [3:0] _GEN_5;
  wire [13:0] _GEN_8;
  wire  _GEN_9;
  wire [31:0] _GEN_10;
  wire [3:0] _GEN_12;
  wire [13:0] _GEN_15;
  wire  _GEN_16;
  wire [31:0] _GEN_17;
  wire [3:0] _GEN_19;
  wire  _T_68;
  wire  _T_69;
  wire  _T_71;
  wire  _T_73;
  wire  _T_75;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  _T_81;
  wire  _T_82;
  assign io_in_1_ready = _T_77;
  assign io_in_2_ready = _T_78;
  assign io_in_3_ready = _T_79;
  assign io_out_valid = _T_82;
  assign io_out_bits_addr = _GEN_15;
  assign io_out_bits_write = _GEN_16;
  assign io_out_bits_wdata = _GEN_17;
  assign io_out_bits_eccMask = _GEN_19;
  assign _GEN_1 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr;
  assign _GEN_2 = io_in_2_valid ? io_in_2_bits_write : io_in_3_bits_write;
  assign _GEN_3 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata;
  assign _GEN_5 = io_in_2_valid ? io_in_2_bits_eccMask : io_in_3_bits_eccMask;
  assign _GEN_8 = io_in_1_valid ? io_in_1_bits_addr : _GEN_1;
  assign _GEN_9 = io_in_1_valid ? io_in_1_bits_write : _GEN_2;
  assign _GEN_10 = io_in_1_valid ? io_in_1_bits_wdata : _GEN_3;
  assign _GEN_12 = io_in_1_valid ? io_in_1_bits_eccMask : _GEN_5;
  assign _GEN_15 = io_in_0_valid ? io_in_0_bits_addr : _GEN_8;
  assign _GEN_16 = io_in_0_valid ? io_in_0_bits_write : _GEN_9;
  assign _GEN_17 = io_in_0_valid ? io_in_0_bits_wdata : _GEN_10;
  assign _GEN_19 = io_in_0_valid ? io_in_0_bits_eccMask : _GEN_12;
  assign _T_68 = io_in_0_valid | io_in_1_valid;
  assign _T_69 = _T_68 | io_in_2_valid;
  assign _T_71 = io_in_0_valid == 1'h0;
  assign _T_73 = _T_68 == 1'h0;
  assign _T_75 = _T_69 == 1'h0;
  assign _T_77 = _T_71 & io_out_ready;
  assign _T_78 = _T_73 & io_out_ready;
  assign _T_79 = _T_75 & io_out_ready;
  assign _T_81 = _T_75 == 1'h0;
  assign _T_82 = _T_81 | io_in_3_valid;
endmodule
module PMPChecker(
  input  [1:0]  io_prv,
  input         io_pmp_0_cfg_l,
  input  [1:0]  io_pmp_0_cfg_a,
  input         io_pmp_0_cfg_x,
  input         io_pmp_0_cfg_w,
  input         io_pmp_0_cfg_r,
  input  [29:0] io_pmp_0_addr,
  input  [31:0] io_pmp_0_mask,
  input         io_pmp_1_cfg_l,
  input  [1:0]  io_pmp_1_cfg_a,
  input         io_pmp_1_cfg_x,
  input         io_pmp_1_cfg_w,
  input         io_pmp_1_cfg_r,
  input  [29:0] io_pmp_1_addr,
  input  [31:0] io_pmp_1_mask,
  input         io_pmp_2_cfg_l,
  input  [1:0]  io_pmp_2_cfg_a,
  input         io_pmp_2_cfg_x,
  input         io_pmp_2_cfg_w,
  input         io_pmp_2_cfg_r,
  input  [29:0] io_pmp_2_addr,
  input  [31:0] io_pmp_2_mask,
  input         io_pmp_3_cfg_l,
  input  [1:0]  io_pmp_3_cfg_a,
  input         io_pmp_3_cfg_x,
  input         io_pmp_3_cfg_w,
  input         io_pmp_3_cfg_r,
  input  [29:0] io_pmp_3_addr,
  input  [31:0] io_pmp_3_mask,
  input         io_pmp_4_cfg_l,
  input  [1:0]  io_pmp_4_cfg_a,
  input         io_pmp_4_cfg_x,
  input         io_pmp_4_cfg_w,
  input         io_pmp_4_cfg_r,
  input  [29:0] io_pmp_4_addr,
  input  [31:0] io_pmp_4_mask,
  input         io_pmp_5_cfg_l,
  input  [1:0]  io_pmp_5_cfg_a,
  input         io_pmp_5_cfg_x,
  input         io_pmp_5_cfg_w,
  input         io_pmp_5_cfg_r,
  input  [29:0] io_pmp_5_addr,
  input  [31:0] io_pmp_5_mask,
  input         io_pmp_6_cfg_l,
  input  [1:0]  io_pmp_6_cfg_a,
  input         io_pmp_6_cfg_x,
  input         io_pmp_6_cfg_w,
  input         io_pmp_6_cfg_r,
  input  [29:0] io_pmp_6_addr,
  input  [31:0] io_pmp_6_mask,
  input         io_pmp_7_cfg_l,
  input  [1:0]  io_pmp_7_cfg_a,
  input         io_pmp_7_cfg_x,
  input         io_pmp_7_cfg_w,
  input         io_pmp_7_cfg_r,
  input  [29:0] io_pmp_7_addr,
  input  [31:0] io_pmp_7_mask,
  input  [31:0] io_addr,
  output        io_r,
  output        io_w,
  output        io_x
);
  wire  default$;
  wire  _T_37;
  wire [31:0] _GEN_0;
  wire [31:0] _T_38;
  wire [31:0] _T_39;
  wire [31:0] _T_40;
  wire [31:0] _T_41;
  wire  _T_43;
  wire  _T_44;
  wire [31:0] _GEN_1;
  wire [31:0] _T_49;
  wire  _T_50;
  wire  _T_52;
  wire  _T_55;
  wire  _T_56;
  wire  _T_57;
  wire  _T_58;
  wire  _T_60;
  wire  _T_61;
  wire  _T_66;
  wire  _T_68;
  wire  _T_70;
  wire  _T_71_cfg_x;
  wire  _T_71_cfg_w;
  wire  _T_71_cfg_r;
  wire  _T_72;
  wire [31:0] _T_74;
  wire [31:0] _T_75;
  wire [31:0] _T_76;
  wire  _T_78;
  wire  _T_79;
  wire [31:0] _GEN_4;
  wire [31:0] _T_84;
  wire  _T_85;
  wire  _T_87;
  wire  _T_91;
  wire  _T_92;
  wire  _T_93;
  wire  _T_95;
  wire  _T_96;
  wire  _T_101;
  wire  _T_103;
  wire  _T_105;
  wire  _T_106_cfg_x;
  wire  _T_106_cfg_w;
  wire  _T_106_cfg_r;
  wire  _T_107;
  wire [31:0] _T_109;
  wire [31:0] _T_110;
  wire [31:0] _T_111;
  wire  _T_113;
  wire  _T_114;
  wire [31:0] _GEN_7;
  wire [31:0] _T_119;
  wire  _T_120;
  wire  _T_122;
  wire  _T_126;
  wire  _T_127;
  wire  _T_128;
  wire  _T_130;
  wire  _T_131;
  wire  _T_136;
  wire  _T_138;
  wire  _T_140;
  wire  _T_141_cfg_x;
  wire  _T_141_cfg_w;
  wire  _T_141_cfg_r;
  wire  _T_142;
  wire [31:0] _T_144;
  wire [31:0] _T_145;
  wire [31:0] _T_146;
  wire  _T_148;
  wire  _T_149;
  wire [31:0] _GEN_10;
  wire [31:0] _T_154;
  wire  _T_155;
  wire  _T_157;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_165;
  wire  _T_166;
  wire  _T_171;
  wire  _T_173;
  wire  _T_175;
  wire  _T_176_cfg_x;
  wire  _T_176_cfg_w;
  wire  _T_176_cfg_r;
  wire  _T_177;
  wire [31:0] _T_179;
  wire [31:0] _T_180;
  wire [31:0] _T_181;
  wire  _T_183;
  wire  _T_184;
  wire [31:0] _GEN_13;
  wire [31:0] _T_189;
  wire  _T_190;
  wire  _T_192;
  wire  _T_196;
  wire  _T_197;
  wire  _T_198;
  wire  _T_200;
  wire  _T_201;
  wire  _T_206;
  wire  _T_208;
  wire  _T_210;
  wire  _T_211_cfg_x;
  wire  _T_211_cfg_w;
  wire  _T_211_cfg_r;
  wire  _T_212;
  wire [31:0] _T_214;
  wire [31:0] _T_215;
  wire [31:0] _T_216;
  wire  _T_218;
  wire  _T_219;
  wire [31:0] _GEN_16;
  wire [31:0] _T_224;
  wire  _T_225;
  wire  _T_227;
  wire  _T_231;
  wire  _T_232;
  wire  _T_233;
  wire  _T_235;
  wire  _T_236;
  wire  _T_241;
  wire  _T_243;
  wire  _T_245;
  wire  _T_246_cfg_x;
  wire  _T_246_cfg_w;
  wire  _T_246_cfg_r;
  wire  _T_247;
  wire [31:0] _T_249;
  wire [31:0] _T_250;
  wire [31:0] _T_251;
  wire  _T_253;
  wire  _T_254;
  wire [31:0] _GEN_19;
  wire [31:0] _T_259;
  wire  _T_260;
  wire  _T_262;
  wire  _T_266;
  wire  _T_267;
  wire  _T_268;
  wire  _T_270;
  wire  _T_271;
  wire  _T_276;
  wire  _T_278;
  wire  _T_280;
  wire  _T_281_cfg_x;
  wire  _T_281_cfg_w;
  wire  _T_281_cfg_r;
  wire  _T_282;
  wire [31:0] _T_284;
  wire [31:0] _T_285;
  wire [31:0] _T_286;
  wire  _T_288;
  wire  _T_289;
  wire  _T_302;
  wire  _T_303;
  wire  _T_305;
  wire  _T_306;
  wire  _T_311;
  wire  _T_313;
  wire  _T_315;
  wire  res_cfg_x;
  wire  res_cfg_w;
  wire  res_cfg_r;
  assign io_r = res_cfg_r;
  assign io_w = res_cfg_w;
  assign io_x = res_cfg_x;
  assign default$ = io_prv > 2'h1;
  assign _T_37 = io_pmp_7_cfg_a[1];
  assign _GEN_0 = {{2'd0}, io_pmp_7_addr};
  assign _T_38 = _GEN_0 << 2;
  assign _T_39 = io_addr ^ _T_38;
  assign _T_40 = ~ io_pmp_7_mask;
  assign _T_41 = _T_39 & _T_40;
  assign _T_43 = _T_41 == 32'h0;
  assign _T_44 = io_pmp_7_cfg_a[0];
  assign _GEN_1 = {{2'd0}, io_pmp_6_addr};
  assign _T_49 = _GEN_1 << 2;
  assign _T_50 = io_addr < _T_49;
  assign _T_52 = _T_50 == 1'h0;
  assign _T_55 = io_addr < _T_38;
  assign _T_56 = _T_52 & _T_55;
  assign _T_57 = _T_44 & _T_56;
  assign _T_58 = _T_37 ? _T_43 : _T_57;
  assign _T_60 = io_pmp_7_cfg_l == 1'h0;
  assign _T_61 = default$ & _T_60;
  assign _T_66 = io_pmp_7_cfg_r | _T_61;
  assign _T_68 = io_pmp_7_cfg_w | _T_61;
  assign _T_70 = io_pmp_7_cfg_x | _T_61;
  assign _T_71_cfg_x = _T_58 ? _T_70 : default$;
  assign _T_71_cfg_w = _T_58 ? _T_68 : default$;
  assign _T_71_cfg_r = _T_58 ? _T_66 : default$;
  assign _T_72 = io_pmp_6_cfg_a[1];
  assign _T_74 = io_addr ^ _T_49;
  assign _T_75 = ~ io_pmp_6_mask;
  assign _T_76 = _T_74 & _T_75;
  assign _T_78 = _T_76 == 32'h0;
  assign _T_79 = io_pmp_6_cfg_a[0];
  assign _GEN_4 = {{2'd0}, io_pmp_5_addr};
  assign _T_84 = _GEN_4 << 2;
  assign _T_85 = io_addr < _T_84;
  assign _T_87 = _T_85 == 1'h0;
  assign _T_91 = _T_87 & _T_50;
  assign _T_92 = _T_79 & _T_91;
  assign _T_93 = _T_72 ? _T_78 : _T_92;
  assign _T_95 = io_pmp_6_cfg_l == 1'h0;
  assign _T_96 = default$ & _T_95;
  assign _T_101 = io_pmp_6_cfg_r | _T_96;
  assign _T_103 = io_pmp_6_cfg_w | _T_96;
  assign _T_105 = io_pmp_6_cfg_x | _T_96;
  assign _T_106_cfg_x = _T_93 ? _T_105 : _T_71_cfg_x;
  assign _T_106_cfg_w = _T_93 ? _T_103 : _T_71_cfg_w;
  assign _T_106_cfg_r = _T_93 ? _T_101 : _T_71_cfg_r;
  assign _T_107 = io_pmp_5_cfg_a[1];
  assign _T_109 = io_addr ^ _T_84;
  assign _T_110 = ~ io_pmp_5_mask;
  assign _T_111 = _T_109 & _T_110;
  assign _T_113 = _T_111 == 32'h0;
  assign _T_114 = io_pmp_5_cfg_a[0];
  assign _GEN_7 = {{2'd0}, io_pmp_4_addr};
  assign _T_119 = _GEN_7 << 2;
  assign _T_120 = io_addr < _T_119;
  assign _T_122 = _T_120 == 1'h0;
  assign _T_126 = _T_122 & _T_85;
  assign _T_127 = _T_114 & _T_126;
  assign _T_128 = _T_107 ? _T_113 : _T_127;
  assign _T_130 = io_pmp_5_cfg_l == 1'h0;
  assign _T_131 = default$ & _T_130;
  assign _T_136 = io_pmp_5_cfg_r | _T_131;
  assign _T_138 = io_pmp_5_cfg_w | _T_131;
  assign _T_140 = io_pmp_5_cfg_x | _T_131;
  assign _T_141_cfg_x = _T_128 ? _T_140 : _T_106_cfg_x;
  assign _T_141_cfg_w = _T_128 ? _T_138 : _T_106_cfg_w;
  assign _T_141_cfg_r = _T_128 ? _T_136 : _T_106_cfg_r;
  assign _T_142 = io_pmp_4_cfg_a[1];
  assign _T_144 = io_addr ^ _T_119;
  assign _T_145 = ~ io_pmp_4_mask;
  assign _T_146 = _T_144 & _T_145;
  assign _T_148 = _T_146 == 32'h0;
  assign _T_149 = io_pmp_4_cfg_a[0];
  assign _GEN_10 = {{2'd0}, io_pmp_3_addr};
  assign _T_154 = _GEN_10 << 2;
  assign _T_155 = io_addr < _T_154;
  assign _T_157 = _T_155 == 1'h0;
  assign _T_161 = _T_157 & _T_120;
  assign _T_162 = _T_149 & _T_161;
  assign _T_163 = _T_142 ? _T_148 : _T_162;
  assign _T_165 = io_pmp_4_cfg_l == 1'h0;
  assign _T_166 = default$ & _T_165;
  assign _T_171 = io_pmp_4_cfg_r | _T_166;
  assign _T_173 = io_pmp_4_cfg_w | _T_166;
  assign _T_175 = io_pmp_4_cfg_x | _T_166;
  assign _T_176_cfg_x = _T_163 ? _T_175 : _T_141_cfg_x;
  assign _T_176_cfg_w = _T_163 ? _T_173 : _T_141_cfg_w;
  assign _T_176_cfg_r = _T_163 ? _T_171 : _T_141_cfg_r;
  assign _T_177 = io_pmp_3_cfg_a[1];
  assign _T_179 = io_addr ^ _T_154;
  assign _T_180 = ~ io_pmp_3_mask;
  assign _T_181 = _T_179 & _T_180;
  assign _T_183 = _T_181 == 32'h0;
  assign _T_184 = io_pmp_3_cfg_a[0];
  assign _GEN_13 = {{2'd0}, io_pmp_2_addr};
  assign _T_189 = _GEN_13 << 2;
  assign _T_190 = io_addr < _T_189;
  assign _T_192 = _T_190 == 1'h0;
  assign _T_196 = _T_192 & _T_155;
  assign _T_197 = _T_184 & _T_196;
  assign _T_198 = _T_177 ? _T_183 : _T_197;
  assign _T_200 = io_pmp_3_cfg_l == 1'h0;
  assign _T_201 = default$ & _T_200;
  assign _T_206 = io_pmp_3_cfg_r | _T_201;
  assign _T_208 = io_pmp_3_cfg_w | _T_201;
  assign _T_210 = io_pmp_3_cfg_x | _T_201;
  assign _T_211_cfg_x = _T_198 ? _T_210 : _T_176_cfg_x;
  assign _T_211_cfg_w = _T_198 ? _T_208 : _T_176_cfg_w;
  assign _T_211_cfg_r = _T_198 ? _T_206 : _T_176_cfg_r;
  assign _T_212 = io_pmp_2_cfg_a[1];
  assign _T_214 = io_addr ^ _T_189;
  assign _T_215 = ~ io_pmp_2_mask;
  assign _T_216 = _T_214 & _T_215;
  assign _T_218 = _T_216 == 32'h0;
  assign _T_219 = io_pmp_2_cfg_a[0];
  assign _GEN_16 = {{2'd0}, io_pmp_1_addr};
  assign _T_224 = _GEN_16 << 2;
  assign _T_225 = io_addr < _T_224;
  assign _T_227 = _T_225 == 1'h0;
  assign _T_231 = _T_227 & _T_190;
  assign _T_232 = _T_219 & _T_231;
  assign _T_233 = _T_212 ? _T_218 : _T_232;
  assign _T_235 = io_pmp_2_cfg_l == 1'h0;
  assign _T_236 = default$ & _T_235;
  assign _T_241 = io_pmp_2_cfg_r | _T_236;
  assign _T_243 = io_pmp_2_cfg_w | _T_236;
  assign _T_245 = io_pmp_2_cfg_x | _T_236;
  assign _T_246_cfg_x = _T_233 ? _T_245 : _T_211_cfg_x;
  assign _T_246_cfg_w = _T_233 ? _T_243 : _T_211_cfg_w;
  assign _T_246_cfg_r = _T_233 ? _T_241 : _T_211_cfg_r;
  assign _T_247 = io_pmp_1_cfg_a[1];
  assign _T_249 = io_addr ^ _T_224;
  assign _T_250 = ~ io_pmp_1_mask;
  assign _T_251 = _T_249 & _T_250;
  assign _T_253 = _T_251 == 32'h0;
  assign _T_254 = io_pmp_1_cfg_a[0];
  assign _GEN_19 = {{2'd0}, io_pmp_0_addr};
  assign _T_259 = _GEN_19 << 2;
  assign _T_260 = io_addr < _T_259;
  assign _T_262 = _T_260 == 1'h0;
  assign _T_266 = _T_262 & _T_225;
  assign _T_267 = _T_254 & _T_266;
  assign _T_268 = _T_247 ? _T_253 : _T_267;
  assign _T_270 = io_pmp_1_cfg_l == 1'h0;
  assign _T_271 = default$ & _T_270;
  assign _T_276 = io_pmp_1_cfg_r | _T_271;
  assign _T_278 = io_pmp_1_cfg_w | _T_271;
  assign _T_280 = io_pmp_1_cfg_x | _T_271;
  assign _T_281_cfg_x = _T_268 ? _T_280 : _T_246_cfg_x;
  assign _T_281_cfg_w = _T_268 ? _T_278 : _T_246_cfg_w;
  assign _T_281_cfg_r = _T_268 ? _T_276 : _T_246_cfg_r;
  assign _T_282 = io_pmp_0_cfg_a[1];
  assign _T_284 = io_addr ^ _T_259;
  assign _T_285 = ~ io_pmp_0_mask;
  assign _T_286 = _T_284 & _T_285;
  assign _T_288 = _T_286 == 32'h0;
  assign _T_289 = io_pmp_0_cfg_a[0];
  assign _T_302 = _T_289 & _T_260;
  assign _T_303 = _T_282 ? _T_288 : _T_302;
  assign _T_305 = io_pmp_0_cfg_l == 1'h0;
  assign _T_306 = default$ & _T_305;
  assign _T_311 = io_pmp_0_cfg_r | _T_306;
  assign _T_313 = io_pmp_0_cfg_w | _T_306;
  assign _T_315 = io_pmp_0_cfg_x | _T_306;
  assign res_cfg_x = _T_303 ? _T_315 : _T_281_cfg_x;
  assign res_cfg_w = _T_303 ? _T_313 : _T_281_cfg_w;
  assign res_cfg_r = _T_303 ? _T_311 : _T_281_cfg_r;
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [31:0] io_req_bits_vaddr,
  input         io_req_bits_instruction,
  input  [1:0]  io_req_bits_size,
  input  [4:0]  io_req_bits_cmd,
  output        io_resp_miss,
  output [31:0] io_resp_paddr,
  output        io_resp_pf_ld,
  output        io_resp_pf_st,
  output        io_resp_pf_inst,
  output        io_resp_ae_ld,
  output        io_resp_ae_st,
  output        io_resp_ae_inst,
  output        io_resp_ma_ld,
  output        io_resp_ma_st,
  output        io_resp_cacheable,
  output        io_ptw_req_valid,
  output [19:0] io_ptw_req_bits_addr,
  input         io_ptw_resp_valid,
  input  [1:0]  io_ptw_status_dprv,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask
);
  reg [53:0] reg_entries_0;
  reg [63:0] _RAND_0;
  reg [53:0] reg_entries_1;
  reg [63:0] _RAND_1;
  reg [53:0] reg_entries_2;
  reg [63:0] _RAND_2;
  reg [53:0] reg_entries_3;
  reg [63:0] _RAND_3;
  reg [53:0] reg_entries_4;
  reg [63:0] _RAND_4;
  wire  _T_68;
  wire  _T_69;
  wire  _T_70;
  wire  _T_71;
  wire  _T_72;
  wire  _T_73;
  wire  _T_74;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_80;
  wire  _T_88;
  wire  _T_89;
  wire  _T_90;
  wire  _T_91;
  wire  _T_92;
  wire  _T_93;
  wire  _T_94;
  wire  _T_95;
  wire  _T_96;
  wire  _T_97;
  wire  _T_100;
  wire  _T_108;
  wire  _T_109;
  wire  _T_110;
  wire  _T_111;
  wire  _T_112;
  wire  _T_113;
  wire  _T_114;
  wire  _T_115;
  wire  _T_116;
  wire  _T_117;
  wire  _T_120;
  wire  _T_128;
  wire  _T_129;
  wire  _T_130;
  wire  _T_131;
  wire  _T_132;
  wire  _T_133;
  wire  _T_134;
  wire  _T_135;
  wire  _T_136;
  wire  _T_137;
  wire  _T_140;
  wire  _T_155;
  wire  _T_156;
  wire  _T_157;
  wire  _T_160;
  reg [1:0] state;
  reg [31:0] _RAND_5;
  reg [19:0] r_refill_tag;
  reg [31:0] _RAND_6;
  wire [1:0] priv;
  wire  priv_s;
  wire [19:0] vpn;
  wire [11:0] pgOffset;
  wire  _T_183;
  wire [31:0] mpu_physaddr;
  wire [1:0] pmp_io_prv;
  wire  pmp_io_pmp_0_cfg_l;
  wire [1:0] pmp_io_pmp_0_cfg_a;
  wire  pmp_io_pmp_0_cfg_x;
  wire  pmp_io_pmp_0_cfg_w;
  wire  pmp_io_pmp_0_cfg_r;
  wire [29:0] pmp_io_pmp_0_addr;
  wire [31:0] pmp_io_pmp_0_mask;
  wire  pmp_io_pmp_1_cfg_l;
  wire [1:0] pmp_io_pmp_1_cfg_a;
  wire  pmp_io_pmp_1_cfg_x;
  wire  pmp_io_pmp_1_cfg_w;
  wire  pmp_io_pmp_1_cfg_r;
  wire [29:0] pmp_io_pmp_1_addr;
  wire [31:0] pmp_io_pmp_1_mask;
  wire  pmp_io_pmp_2_cfg_l;
  wire [1:0] pmp_io_pmp_2_cfg_a;
  wire  pmp_io_pmp_2_cfg_x;
  wire  pmp_io_pmp_2_cfg_w;
  wire  pmp_io_pmp_2_cfg_r;
  wire [29:0] pmp_io_pmp_2_addr;
  wire [31:0] pmp_io_pmp_2_mask;
  wire  pmp_io_pmp_3_cfg_l;
  wire [1:0] pmp_io_pmp_3_cfg_a;
  wire  pmp_io_pmp_3_cfg_x;
  wire  pmp_io_pmp_3_cfg_w;
  wire  pmp_io_pmp_3_cfg_r;
  wire [29:0] pmp_io_pmp_3_addr;
  wire [31:0] pmp_io_pmp_3_mask;
  wire  pmp_io_pmp_4_cfg_l;
  wire [1:0] pmp_io_pmp_4_cfg_a;
  wire  pmp_io_pmp_4_cfg_x;
  wire  pmp_io_pmp_4_cfg_w;
  wire  pmp_io_pmp_4_cfg_r;
  wire [29:0] pmp_io_pmp_4_addr;
  wire [31:0] pmp_io_pmp_4_mask;
  wire  pmp_io_pmp_5_cfg_l;
  wire [1:0] pmp_io_pmp_5_cfg_a;
  wire  pmp_io_pmp_5_cfg_x;
  wire  pmp_io_pmp_5_cfg_w;
  wire  pmp_io_pmp_5_cfg_r;
  wire [29:0] pmp_io_pmp_5_addr;
  wire [31:0] pmp_io_pmp_5_mask;
  wire  pmp_io_pmp_6_cfg_l;
  wire [1:0] pmp_io_pmp_6_cfg_a;
  wire  pmp_io_pmp_6_cfg_x;
  wire  pmp_io_pmp_6_cfg_w;
  wire  pmp_io_pmp_6_cfg_r;
  wire [29:0] pmp_io_pmp_6_addr;
  wire [31:0] pmp_io_pmp_6_mask;
  wire  pmp_io_pmp_7_cfg_l;
  wire [1:0] pmp_io_pmp_7_cfg_a;
  wire  pmp_io_pmp_7_cfg_x;
  wire  pmp_io_pmp_7_cfg_w;
  wire  pmp_io_pmp_7_cfg_r;
  wire [29:0] pmp_io_pmp_7_addr;
  wire [31:0] pmp_io_pmp_7_mask;
  wire [31:0] pmp_io_addr;
  wire  pmp_io_r;
  wire  pmp_io_w;
  wire  pmp_io_x;
  wire [31:0] _T_193;
  wire [32:0] _T_194;
  wire [32:0] _T_196;
  wire [32:0] _T_197;
  wire  _T_199;
  wire [31:0] _T_201;
  wire [32:0] _T_202;
  wire [32:0] _T_204;
  wire [32:0] _T_205;
  wire  _T_207;
  wire [32:0] _T_210;
  wire [32:0] _T_212;
  wire [32:0] _T_213;
  wire  _T_215;
  wire [31:0] _T_217;
  wire [32:0] _T_218;
  wire [32:0] _T_220;
  wire [32:0] _T_221;
  wire  _T_223;
  wire [31:0] _T_225;
  wire [32:0] _T_226;
  wire [32:0] _T_228;
  wire [32:0] _T_229;
  wire  _T_231;
  wire [31:0] _T_233;
  wire [32:0] _T_234;
  wire [32:0] _T_236;
  wire [32:0] _T_237;
  wire  _T_239;
  wire [31:0] _T_241;
  wire [32:0] _T_242;
  wire [32:0] _T_244;
  wire [32:0] _T_245;
  wire  _T_247;
  wire  _T_260;
  wire  _T_261;
  wire  _T_262;
  wire  _T_263;
  wire  _T_264;
  wire  legal_address;
  wire [32:0] _T_269;
  wire [32:0] _T_270;
  wire  _T_272;
  wire [32:0] _T_277;
  wire [32:0] _T_278;
  wire  _T_280;
  wire [32:0] _T_285;
  wire [32:0] _T_286;
  wire  _T_288;
  wire [32:0] _T_293;
  wire [32:0] _T_294;
  wire  _T_296;
  wire [32:0] _T_301;
  wire [32:0] _T_302;
  wire  _T_304;
  wire [32:0] _T_309;
  wire [32:0] _T_310;
  wire  _T_312;
  wire  _T_313;
  wire  _T_314;
  wire [31:0] _T_320;
  wire [32:0] _T_321;
  wire [32:0] _T_323;
  wire [32:0] _T_324;
  wire  _T_326;
  wire  cacheable;
  wire  prot_r;
  wire [31:0] _T_356;
  wire [32:0] _T_357;
  wire [32:0] _T_359;
  wire [32:0] _T_360;
  wire  _T_362;
  wire [32:0] _T_367;
  wire [32:0] _T_368;
  wire  _T_370;
  wire [32:0] _T_375;
  wire [32:0] _T_376;
  wire  _T_378;
  wire  _T_379;
  wire  _T_380;
  wire  _T_390;
  wire  prot_w;
  wire  _T_435;
  wire  prot_al;
  wire  _T_540;
  wire  _T_541;
  wire  _T_542;
  wire  _T_552;
  wire  prot_x;
  wire  _T_614;
  wire  prot_eff;
  wire [9:0] _T_629;
  wire [9:0] _T_636;
  wire [19:0] ppn;
  wire  _T_836;
  wire  _T_837;
  wire [1:0] _T_838;
  wire [1:0] _T_839;
  wire [2:0] _T_840;
  wire [4:0] _T_841;
  wire [4:0] _T_843;
  wire [4:0] _T_848;
  wire [4:0] _T_850;
  wire [4:0] priv_rw_ok;
  wire [4:0] priv_x_ok;
  wire [1:0] _T_861;
  wire [1:0] _T_862;
  wire [2:0] _T_863;
  wire [4:0] _T_864;
  wire [1:0] _T_865;
  wire [1:0] _T_866;
  wire [2:0] _T_867;
  wire [4:0] _T_868;
  wire [4:0] _T_870;
  wire [4:0] _T_871;
  wire [4:0] _T_872;
  wire [5:0] r_array;
  wire [1:0] _T_874;
  wire [1:0] _T_875;
  wire [2:0] _T_876;
  wire [4:0] _T_877;
  wire [4:0] _T_878;
  wire [5:0] w_array;
  wire [4:0] _T_884;
  wire [5:0] x_array;
  wire [1:0] _T_888;
  wire [1:0] _T_889;
  wire [1:0] _T_890;
  wire [3:0] _T_891;
  wire [5:0] pr_array;
  wire [1:0] _T_895;
  wire [1:0] _T_896;
  wire [1:0] _T_897;
  wire [3:0] _T_898;
  wire [5:0] pw_array;
  wire [1:0] _T_902;
  wire [1:0] _T_903;
  wire [1:0] _T_904;
  wire [3:0] _T_905;
  wire [5:0] px_array;
  wire [1:0] _T_909;
  wire [1:0] _T_910;
  wire [1:0] _T_911;
  wire [3:0] _T_912;
  wire [5:0] paa_array;
  wire [1:0] _T_917;
  wire [1:0] _T_918;
  wire [3:0] _T_919;
  wire [5:0] pal_array;
  wire [1:0] _T_923;
  wire [1:0] _T_924;
  wire [1:0] _T_925;
  wire [3:0] _T_926;
  wire [5:0] eff_array;
  wire [1:0] _T_930;
  wire [1:0] _T_931;
  wire [1:0] _T_932;
  wire [3:0] _T_933;
  wire [5:0] c_array;
  wire [3:0] _T_935;
  wire [4:0] _T_937;
  wire [4:0] _T_938;
  wire [3:0] _T_939;
  wire [31:0] _GEN_14;
  wire [31:0] _T_940;
  wire  misaligned;
  wire [5:0] _T_946;
  wire  _T_950;
  wire  _T_951;
  wire  _T_952;
  wire [5:0] _T_956;
  wire [5:0] ae_array;
  wire  _T_958;
  wire  _T_961;
  wire  _T_964;
  wire  _T_969;
  wire  _T_970;
  wire  _T_971;
  wire  _T_972;
  wire  _T_973;
  wire  _T_974;
  wire  _T_975;
  wire  _T_981;
  wire  _T_982;
  wire  _T_983;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire  _T_987;
  wire  _T_988;
  wire  _T_989;
  wire  _T_990;
  wire  _T_991;
  wire [5:0] _T_992;
  wire [5:0] _T_993;
  wire [5:0] ae_ld_array;
  wire  _T_996;
  wire  _T_998;
  wire  _T_999;
  wire  _T_1002;
  wire  _T_1029;
  wire [5:0] _T_1030;
  wire [5:0] _T_1031;
  wire [5:0] _T_1033;
  wire [5:0] _T_1047;
  wire [5:0] _T_1049;
  wire [5:0] _T_1050;
  wire [5:0] _T_1067;
  wire [5:0] _T_1069;
  wire [5:0] ae_st_array;
  wire  _T_1105;
  wire [5:0] _T_1106;
  wire [5:0] ma_ld_array;
  wire  _T_1143;
  wire [5:0] ma_st_array;
  wire [5:0] _GEN_15;
  wire [5:0] _T_1181;
  wire [5:0] _T_1182;
  wire [5:0] pf_ld_array;
  wire [5:0] _T_1219;
  wire [5:0] _T_1220;
  wire [5:0] pf_st_array;
  wire [5:0] _T_1222;
  wire [5:0] pf_inst_array;
  wire  _T_1305;
  wire [5:0] _T_1342;
  wire  _T_1344;
  wire [5:0] _T_1382;
  wire  _T_1384;
  wire [5:0] _T_1386;
  wire  _T_1388;
  wire [5:0] _T_1390;
  wire  _T_1392;
  wire [5:0] _T_1393;
  wire  _T_1395;
  wire [5:0] _T_1396;
  wire [5:0] _T_1397;
  wire  _T_1399;
  wire [5:0] _T_1400;
  wire  _T_1402;
  wire [5:0] _T_1403;
  wire  _T_1405;
  wire [5:0] _T_1407;
  wire  _T_1409;
  wire [31:0] _T_1412;
  PMPChecker pmp (
    .io_prv(pmp_io_prv),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_addr(pmp_io_addr),
    .io_r(pmp_io_r),
    .io_w(pmp_io_w),
    .io_x(pmp_io_x)
  );
  assign io_req_ready = _T_1305;
  assign io_resp_miss = 1'h0;
  assign io_resp_paddr = _T_1412;
  assign io_resp_pf_ld = _T_1344;
  assign io_resp_pf_st = _T_1384;
  assign io_resp_pf_inst = _T_1388;
  assign io_resp_ae_ld = _T_1392;
  assign io_resp_ae_st = _T_1395;
  assign io_resp_ae_inst = _T_1399;
  assign io_resp_ma_ld = _T_1402;
  assign io_resp_ma_st = _T_1405;
  assign io_resp_cacheable = _T_1409;
  assign io_ptw_req_valid = _T_183;
  assign io_ptw_req_bits_addr = r_refill_tag;
  assign _T_68 = reg_entries_0[0];
  assign _T_69 = reg_entries_0[1];
  assign _T_70 = reg_entries_0[2];
  assign _T_71 = reg_entries_0[3];
  assign _T_72 = reg_entries_0[4];
  assign _T_73 = reg_entries_0[5];
  assign _T_74 = reg_entries_0[6];
  assign _T_75 = reg_entries_0[7];
  assign _T_76 = reg_entries_0[8];
  assign _T_77 = reg_entries_0[9];
  assign _T_78 = reg_entries_0[10];
  assign _T_80 = reg_entries_0[12];
  assign _T_88 = reg_entries_1[0];
  assign _T_89 = reg_entries_1[1];
  assign _T_90 = reg_entries_1[2];
  assign _T_91 = reg_entries_1[3];
  assign _T_92 = reg_entries_1[4];
  assign _T_93 = reg_entries_1[5];
  assign _T_94 = reg_entries_1[6];
  assign _T_95 = reg_entries_1[7];
  assign _T_96 = reg_entries_1[8];
  assign _T_97 = reg_entries_1[9];
  assign _T_100 = reg_entries_1[12];
  assign _T_108 = reg_entries_2[0];
  assign _T_109 = reg_entries_2[1];
  assign _T_110 = reg_entries_2[2];
  assign _T_111 = reg_entries_2[3];
  assign _T_112 = reg_entries_2[4];
  assign _T_113 = reg_entries_2[5];
  assign _T_114 = reg_entries_2[6];
  assign _T_115 = reg_entries_2[7];
  assign _T_116 = reg_entries_2[8];
  assign _T_117 = reg_entries_2[9];
  assign _T_120 = reg_entries_2[12];
  assign _T_128 = reg_entries_3[0];
  assign _T_129 = reg_entries_3[1];
  assign _T_130 = reg_entries_3[2];
  assign _T_131 = reg_entries_3[3];
  assign _T_132 = reg_entries_3[4];
  assign _T_133 = reg_entries_3[5];
  assign _T_134 = reg_entries_3[6];
  assign _T_135 = reg_entries_3[7];
  assign _T_136 = reg_entries_3[8];
  assign _T_137 = reg_entries_3[9];
  assign _T_140 = reg_entries_3[12];
  assign _T_155 = reg_entries_4[7];
  assign _T_156 = reg_entries_4[8];
  assign _T_157 = reg_entries_4[9];
  assign _T_160 = reg_entries_4[12];
  assign priv = io_req_bits_instruction ? io_ptw_status_prv : io_ptw_status_dprv;
  assign priv_s = priv[0];
  assign vpn = io_req_bits_vaddr[31:12];
  assign pgOffset = io_req_bits_vaddr[11:0];
  assign _T_183 = state == 2'h1;
  assign mpu_physaddr = {vpn,pgOffset};
  assign pmp_io_prv = priv;
  assign pmp_io_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
  assign pmp_io_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
  assign pmp_io_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
  assign pmp_io_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
  assign pmp_io_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
  assign pmp_io_pmp_0_addr = io_ptw_pmp_0_addr;
  assign pmp_io_pmp_0_mask = io_ptw_pmp_0_mask;
  assign pmp_io_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
  assign pmp_io_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
  assign pmp_io_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
  assign pmp_io_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
  assign pmp_io_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
  assign pmp_io_pmp_1_addr = io_ptw_pmp_1_addr;
  assign pmp_io_pmp_1_mask = io_ptw_pmp_1_mask;
  assign pmp_io_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
  assign pmp_io_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
  assign pmp_io_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
  assign pmp_io_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
  assign pmp_io_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
  assign pmp_io_pmp_2_addr = io_ptw_pmp_2_addr;
  assign pmp_io_pmp_2_mask = io_ptw_pmp_2_mask;
  assign pmp_io_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
  assign pmp_io_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
  assign pmp_io_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
  assign pmp_io_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
  assign pmp_io_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
  assign pmp_io_pmp_3_addr = io_ptw_pmp_3_addr;
  assign pmp_io_pmp_3_mask = io_ptw_pmp_3_mask;
  assign pmp_io_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
  assign pmp_io_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
  assign pmp_io_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
  assign pmp_io_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
  assign pmp_io_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
  assign pmp_io_pmp_4_addr = io_ptw_pmp_4_addr;
  assign pmp_io_pmp_4_mask = io_ptw_pmp_4_mask;
  assign pmp_io_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
  assign pmp_io_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
  assign pmp_io_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
  assign pmp_io_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
  assign pmp_io_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
  assign pmp_io_pmp_5_addr = io_ptw_pmp_5_addr;
  assign pmp_io_pmp_5_mask = io_ptw_pmp_5_mask;
  assign pmp_io_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
  assign pmp_io_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
  assign pmp_io_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
  assign pmp_io_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
  assign pmp_io_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
  assign pmp_io_pmp_6_addr = io_ptw_pmp_6_addr;
  assign pmp_io_pmp_6_mask = io_ptw_pmp_6_mask;
  assign pmp_io_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
  assign pmp_io_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
  assign pmp_io_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
  assign pmp_io_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
  assign pmp_io_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
  assign pmp_io_pmp_7_addr = io_ptw_pmp_7_addr;
  assign pmp_io_pmp_7_mask = io_ptw_pmp_7_mask;
  assign pmp_io_addr = mpu_physaddr;
  assign _T_193 = mpu_physaddr ^ 32'hc000000;
  assign _T_194 = {1'b0,$signed(_T_193)};
  assign _T_196 = $signed(_T_194) & $signed(-33'sh4000000);
  assign _T_197 = $signed(_T_196);
  assign _T_199 = $signed(_T_197) == $signed(33'sh0);
  assign _T_201 = mpu_physaddr ^ 32'h2000000;
  assign _T_202 = {1'b0,$signed(_T_201)};
  assign _T_204 = $signed(_T_202) & $signed(-33'sh10000);
  assign _T_205 = $signed(_T_204);
  assign _T_207 = $signed(_T_205) == $signed(33'sh0);
  assign _T_210 = {1'b0,$signed(mpu_physaddr)};
  assign _T_212 = $signed(_T_210) & $signed(-33'sh1000);
  assign _T_213 = $signed(_T_212);
  assign _T_215 = $signed(_T_213) == $signed(33'sh0);
  assign _T_217 = mpu_physaddr ^ 32'h10000;
  assign _T_218 = {1'b0,$signed(_T_217)};
  assign _T_220 = $signed(_T_218) & $signed(-33'sh10000);
  assign _T_221 = $signed(_T_220);
  assign _T_223 = $signed(_T_221) == $signed(33'sh0);
  assign _T_225 = mpu_physaddr ^ 32'h80000000;
  assign _T_226 = {1'b0,$signed(_T_225)};
  assign _T_228 = $signed(_T_226) & $signed(-33'sh4000);
  assign _T_229 = $signed(_T_228);
  assign _T_231 = $signed(_T_229) == $signed(33'sh0);
  assign _T_233 = mpu_physaddr ^ 32'h60000000;
  assign _T_234 = {1'b0,$signed(_T_233)};
  assign _T_236 = $signed(_T_234) & $signed(-33'sh20000000);
  assign _T_237 = $signed(_T_236);
  assign _T_239 = $signed(_T_237) == $signed(33'sh0);
  assign _T_241 = mpu_physaddr ^ 32'h3000;
  assign _T_242 = {1'b0,$signed(_T_241)};
  assign _T_244 = $signed(_T_242) & $signed(-33'sh1000);
  assign _T_245 = $signed(_T_244);
  assign _T_247 = $signed(_T_245) == $signed(33'sh0);
  assign _T_260 = _T_199 | _T_207;
  assign _T_261 = _T_260 | _T_215;
  assign _T_262 = _T_261 | _T_223;
  assign _T_263 = _T_262 | _T_231;
  assign _T_264 = _T_263 | _T_239;
  assign legal_address = _T_264 | _T_247;
  assign _T_269 = $signed(_T_194) & $signed(33'shfc000000);
  assign _T_270 = $signed(_T_269);
  assign _T_272 = $signed(_T_270) == $signed(33'sh0);
  assign _T_277 = $signed(_T_202) & $signed(33'shffff0000);
  assign _T_278 = $signed(_T_277);
  assign _T_280 = $signed(_T_278) == $signed(33'sh0);
  assign _T_285 = $signed(_T_210) & $signed(33'shffffd000);
  assign _T_286 = $signed(_T_285);
  assign _T_288 = $signed(_T_286) == $signed(33'sh0);
  assign _T_293 = $signed(_T_218) & $signed(33'shffff0000);
  assign _T_294 = $signed(_T_293);
  assign _T_296 = $signed(_T_294) == $signed(33'sh0);
  assign _T_301 = $signed(_T_226) & $signed(33'shffffc000);
  assign _T_302 = $signed(_T_301);
  assign _T_304 = $signed(_T_302) == $signed(33'sh0);
  assign _T_309 = $signed(_T_234) & $signed(33'she0000000);
  assign _T_310 = $signed(_T_309);
  assign _T_312 = $signed(_T_310) == $signed(33'sh0);
  assign _T_313 = _T_272 | _T_280;
  assign _T_314 = _T_313 | _T_288;
  assign _T_320 = mpu_physaddr ^ 32'h1000;
  assign _T_321 = {1'b0,$signed(_T_320)};
  assign _T_323 = $signed(_T_321) & $signed(33'shffffd000);
  assign _T_324 = $signed(_T_323);
  assign _T_326 = $signed(_T_324) == $signed(33'sh0);
  assign cacheable = legal_address & _T_326;
  assign prot_r = legal_address & pmp_io_r;
  assign _T_356 = mpu_physaddr ^ 32'h4000000;
  assign _T_357 = {1'b0,$signed(_T_356)};
  assign _T_359 = $signed(_T_357) & $signed(33'sh74000000);
  assign _T_360 = $signed(_T_359);
  assign _T_362 = $signed(_T_360) == $signed(33'sh0);
  assign _T_367 = $signed(_T_210) & $signed(33'sh74010000);
  assign _T_368 = $signed(_T_367);
  assign _T_370 = $signed(_T_368) == $signed(33'sh0);
  assign _T_375 = $signed(_T_234) & $signed(33'sh60000000);
  assign _T_376 = $signed(_T_375);
  assign _T_378 = $signed(_T_376) == $signed(33'sh0);
  assign _T_379 = _T_362 | _T_370;
  assign _T_380 = _T_379 | _T_378;
  assign _T_390 = legal_address & _T_380;
  assign prot_w = _T_390 & pmp_io_w;
  assign _T_435 = legal_address & _T_379;
  assign prot_al = _T_435 | cacheable;
  assign _T_540 = _T_288 | _T_296;
  assign _T_541 = _T_540 | _T_304;
  assign _T_542 = _T_541 | _T_312;
  assign _T_552 = legal_address & _T_542;
  assign prot_x = _T_552 & pmp_io_x;
  assign _T_614 = _T_314 | _T_312;
  assign prot_eff = legal_address & _T_614;
  assign _T_629 = vpn[19:10];
  assign _T_636 = vpn[9:0];
  assign ppn = {_T_629,_T_636};
  assign _T_836 = priv_s == 1'h0;
  assign _T_837 = _T_836 | io_ptw_status_sum;
  assign _T_838 = {_T_100,_T_80};
  assign _T_839 = {_T_160,_T_140};
  assign _T_840 = {_T_839,_T_120};
  assign _T_841 = {_T_840,_T_838};
  assign _T_843 = _T_837 ? _T_841 : 5'h0;
  assign _T_848 = ~ _T_841;
  assign _T_850 = priv_s ? _T_848 : 5'h0;
  assign priv_rw_ok = _T_843 | _T_850;
  assign priv_x_ok = priv_s ? _T_848 : _T_841;
  assign _T_861 = {_T_95,_T_75};
  assign _T_862 = {_T_155,_T_135};
  assign _T_863 = {_T_862,_T_115};
  assign _T_864 = {_T_863,_T_861};
  assign _T_865 = {_T_96,_T_76};
  assign _T_866 = {_T_156,_T_136};
  assign _T_867 = {_T_866,_T_116};
  assign _T_868 = {_T_867,_T_865};
  assign _T_870 = io_ptw_status_mxr ? _T_868 : 5'h0;
  assign _T_871 = _T_864 | _T_870;
  assign _T_872 = priv_rw_ok & _T_871;
  assign r_array = {1'h1,_T_872};
  assign _T_874 = {_T_97,_T_77};
  assign _T_875 = {_T_157,_T_137};
  assign _T_876 = {_T_875,_T_117};
  assign _T_877 = {_T_876,_T_874};
  assign _T_878 = priv_rw_ok & _T_877;
  assign w_array = {1'h1,_T_878};
  assign _T_884 = priv_x_ok & _T_868;
  assign x_array = {1'h1,_T_884};
  assign _T_888 = prot_r ? 2'h3 : 2'h0;
  assign _T_889 = {_T_92,_T_72};
  assign _T_890 = {_T_132,_T_112};
  assign _T_891 = {_T_890,_T_889};
  assign pr_array = {_T_888,_T_891};
  assign _T_895 = prot_w ? 2'h3 : 2'h0;
  assign _T_896 = {_T_94,_T_74};
  assign _T_897 = {_T_134,_T_114};
  assign _T_898 = {_T_897,_T_896};
  assign pw_array = {_T_895,_T_898};
  assign _T_902 = prot_x ? 2'h3 : 2'h0;
  assign _T_903 = {_T_93,_T_73};
  assign _T_904 = {_T_133,_T_113};
  assign _T_905 = {_T_904,_T_903};
  assign px_array = {_T_902,_T_905};
  assign _T_909 = prot_al ? 2'h3 : 2'h0;
  assign _T_910 = {_T_90,_T_70};
  assign _T_911 = {_T_130,_T_110};
  assign _T_912 = {_T_911,_T_910};
  assign paa_array = {_T_909,_T_912};
  assign _T_917 = {_T_91,_T_71};
  assign _T_918 = {_T_131,_T_111};
  assign _T_919 = {_T_918,_T_917};
  assign pal_array = {_T_909,_T_919};
  assign _T_923 = prot_eff ? 2'h3 : 2'h0;
  assign _T_924 = {_T_89,_T_69};
  assign _T_925 = {_T_129,_T_109};
  assign _T_926 = {_T_925,_T_924};
  assign eff_array = {_T_923,_T_926};
  assign _T_930 = cacheable ? 2'h3 : 2'h0;
  assign _T_931 = {_T_88,_T_68};
  assign _T_932 = {_T_128,_T_108};
  assign _T_933 = {_T_932,_T_931};
  assign c_array = {_T_930,_T_933};
  assign _T_935 = 4'h1 << io_req_bits_size;
  assign _T_937 = _T_935 - 4'h1;
  assign _T_938 = $unsigned(_T_937);
  assign _T_939 = _T_938[3:0];
  assign _GEN_14 = {{28'd0}, _T_939};
  assign _T_940 = io_req_bits_vaddr & _GEN_14;
  assign misaligned = _T_940 != 32'h0;
  assign _T_946 = misaligned ? eff_array : 6'h0;
  assign _T_950 = io_req_bits_cmd == 5'h6;
  assign _T_951 = io_req_bits_cmd == 5'h7;
  assign _T_952 = _T_950 | _T_951;
  assign _T_956 = _T_952 ? 6'h3f : 6'h0;
  assign ae_array = _T_946 | _T_956;
  assign _T_958 = io_req_bits_cmd == 5'h0;
  assign _T_961 = _T_958 | _T_950;
  assign _T_964 = _T_961 | _T_951;
  assign _T_969 = io_req_bits_cmd == 5'h4;
  assign _T_970 = io_req_bits_cmd == 5'h9;
  assign _T_971 = io_req_bits_cmd == 5'ha;
  assign _T_972 = io_req_bits_cmd == 5'hb;
  assign _T_973 = _T_969 | _T_970;
  assign _T_974 = _T_973 | _T_971;
  assign _T_975 = _T_974 | _T_972;
  assign _T_981 = io_req_bits_cmd == 5'h8;
  assign _T_982 = io_req_bits_cmd == 5'hc;
  assign _T_983 = io_req_bits_cmd == 5'hd;
  assign _T_984 = io_req_bits_cmd == 5'he;
  assign _T_985 = io_req_bits_cmd == 5'hf;
  assign _T_986 = _T_981 | _T_982;
  assign _T_987 = _T_986 | _T_983;
  assign _T_988 = _T_987 | _T_984;
  assign _T_989 = _T_988 | _T_985;
  assign _T_990 = _T_975 | _T_989;
  assign _T_991 = _T_964 | _T_990;
  assign _T_992 = ~ pr_array;
  assign _T_993 = ae_array | _T_992;
  assign ae_ld_array = _T_991 ? _T_993 : 6'h0;
  assign _T_996 = io_req_bits_cmd == 5'h1;
  assign _T_998 = io_req_bits_cmd == 5'h11;
  assign _T_999 = _T_996 | _T_998;
  assign _T_1002 = _T_999 | _T_951;
  assign _T_1029 = _T_1002 | _T_990;
  assign _T_1030 = ~ pw_array;
  assign _T_1031 = ae_array | _T_1030;
  assign _T_1033 = _T_1029 ? _T_1031 : 6'h0;
  assign _T_1047 = ~ pal_array;
  assign _T_1049 = _T_975 ? _T_1047 : 6'h0;
  assign _T_1050 = _T_1033 | _T_1049;
  assign _T_1067 = ~ paa_array;
  assign _T_1069 = _T_989 ? _T_1067 : 6'h0;
  assign ae_st_array = _T_1050 | _T_1069;
  assign _T_1105 = misaligned & _T_991;
  assign _T_1106 = ~ eff_array;
  assign ma_ld_array = _T_1105 ? _T_1106 : 6'h0;
  assign _T_1143 = misaligned & _T_1029;
  assign ma_st_array = _T_1143 ? _T_1106 : 6'h0;
  assign _GEN_15 = {{5'd0}, _T_78};
  assign _T_1181 = r_array | _GEN_15;
  assign _T_1182 = ~ _T_1181;
  assign pf_ld_array = _T_991 ? _T_1182 : 6'h0;
  assign _T_1219 = w_array | _GEN_15;
  assign _T_1220 = ~ _T_1219;
  assign pf_st_array = _T_1029 ? _T_1220 : 6'h0;
  assign _T_1222 = x_array | _GEN_15;
  assign pf_inst_array = ~ _T_1222;
  assign _T_1305 = state == 2'h0;
  assign _T_1342 = pf_ld_array & 6'h20;
  assign _T_1344 = _T_1342 != 6'h0;
  assign _T_1382 = pf_st_array & 6'h20;
  assign _T_1384 = _T_1382 != 6'h0;
  assign _T_1386 = pf_inst_array & 6'h20;
  assign _T_1388 = _T_1386 != 6'h0;
  assign _T_1390 = ae_ld_array & 6'h20;
  assign _T_1392 = _T_1390 != 6'h0;
  assign _T_1393 = ae_st_array & 6'h20;
  assign _T_1395 = _T_1393 != 6'h0;
  assign _T_1396 = ~ px_array;
  assign _T_1397 = _T_1396 & 6'h20;
  assign _T_1399 = _T_1397 != 6'h0;
  assign _T_1400 = ma_ld_array & 6'h20;
  assign _T_1402 = _T_1400 != 6'h0;
  assign _T_1403 = ma_st_array & 6'h20;
  assign _T_1405 = _T_1403 != 6'h0;
  assign _T_1407 = c_array & 6'h20;
  assign _T_1409 = _T_1407 != 6'h0;
  assign _T_1412 = {ppn,pgOffset};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{$random}};
  reg_entries_0 = _RAND_0[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{$random}};
  reg_entries_1 = _RAND_1[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{$random}};
  reg_entries_2 = _RAND_2[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{$random}};
  reg_entries_3 = _RAND_3[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{$random}};
  reg_entries_4 = _RAND_4[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  state = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  r_refill_tag = _RAND_6[19:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end
  end
endmodule
module AMOALU(
  input  [3:0]  io_mask,
  input  [4:0]  io_cmd,
  input  [31:0] io_lhs,
  input  [31:0] io_rhs,
  output [31:0] io_out
);
  wire  _T_8;
  wire  _T_10;
  wire  max;
  wire  _T_12;
  wire  _T_14;
  wire  min;
  wire  add;
  wire  _T_17;
  wire  _T_19;
  wire  logic_and;
  wire  _T_21;
  wire  logic_xor;
  wire [32:0] _T_24;
  wire [31:0] adder_out;
  wire [4:0] _T_28;
  wire  _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_34;
  wire  _T_35;
  wire  _T_38;
  wire  less;
  wire  _T_39;
  wire [31:0] minmax;
  wire [31:0] _T_40;
  wire [31:0] _T_42;
  wire [31:0] _T_43;
  wire [31:0] _T_45;
  wire [31:0] logic$;
  wire  _T_46;
  wire [31:0] _T_47;
  wire [31:0] out;
  wire  _T_48;
  wire  _T_49;
  wire  _T_50;
  wire  _T_51;
  wire [7:0] _T_55;
  wire [7:0] _T_59;
  wire [7:0] _T_63;
  wire [7:0] _T_67;
  wire [15:0] _T_68;
  wire [15:0] _T_69;
  wire [31:0] wmask;
  wire [31:0] _T_70;
  wire [31:0] _T_71;
  wire [31:0] _T_72;
  wire [31:0] _T_73;
  assign io_out = _T_73;
  assign _T_8 = io_cmd == 5'hd;
  assign _T_10 = io_cmd == 5'hf;
  assign max = _T_8 | _T_10;
  assign _T_12 = io_cmd == 5'hc;
  assign _T_14 = io_cmd == 5'he;
  assign min = _T_12 | _T_14;
  assign add = io_cmd == 5'h8;
  assign _T_17 = io_cmd == 5'ha;
  assign _T_19 = io_cmd == 5'hb;
  assign logic_and = _T_17 | _T_19;
  assign _T_21 = io_cmd == 5'h9;
  assign logic_xor = _T_21 | _T_17;
  assign _T_24 = io_lhs + io_rhs;
  assign adder_out = _T_24[31:0];
  assign _T_28 = io_cmd & 5'h2;
  assign _T_31 = _T_28 == 5'h0;
  assign _T_32 = io_lhs[31];
  assign _T_33 = io_rhs[31];
  assign _T_34 = _T_32 == _T_33;
  assign _T_35 = io_lhs < io_rhs;
  assign _T_38 = _T_31 ? _T_32 : _T_33;
  assign less = _T_34 ? _T_35 : _T_38;
  assign _T_39 = less ? min : max;
  assign minmax = _T_39 ? io_lhs : io_rhs;
  assign _T_40 = io_lhs & io_rhs;
  assign _T_42 = logic_and ? _T_40 : 32'h0;
  assign _T_43 = io_lhs ^ io_rhs;
  assign _T_45 = logic_xor ? _T_43 : 32'h0;
  assign logic$ = _T_42 | _T_45;
  assign _T_46 = logic_and | logic_xor;
  assign _T_47 = _T_46 ? logic$ : minmax;
  assign out = add ? adder_out : _T_47;
  assign _T_48 = io_mask[0];
  assign _T_49 = io_mask[1];
  assign _T_50 = io_mask[2];
  assign _T_51 = io_mask[3];
  assign _T_55 = _T_48 ? 8'hff : 8'h0;
  assign _T_59 = _T_49 ? 8'hff : 8'h0;
  assign _T_63 = _T_50 ? 8'hff : 8'h0;
  assign _T_67 = _T_51 ? 8'hff : 8'h0;
  assign _T_68 = {_T_59,_T_55};
  assign _T_69 = {_T_67,_T_63};
  assign wmask = {_T_69,_T_68};
  assign _T_70 = wmask & out;
  assign _T_71 = ~ wmask;
  assign _T_72 = _T_71 & io_lhs;
  assign _T_73 = _T_70 | _T_72;
endmodule
module DCache_dcache(
  input         clock,
  input         reset,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [6:0]  io_cpu_req_bits_tag,
  input  [4:0]  io_cpu_req_bits_cmd,
  input  [2:0]  io_cpu_req_bits_typ,
  input         io_cpu_req_bits_phys,
  input         io_cpu_s1_kill,
  input  [31:0] io_cpu_s1_data_data,
  input  [3:0]  io_cpu_s1_data_mask,
  output        io_cpu_s2_nack,
  output        io_cpu_resp_valid,
  output [6:0]  io_cpu_resp_bits_tag,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_replay,
  output        io_cpu_resp_bits_has_data,
  output [31:0] io_cpu_resp_bits_data_word_bypass,
  output [31:0] io_cpu_resp_bits_data_raw,
  output        io_cpu_replay_next,
  output        io_cpu_s2_xcpt_ma_ld,
  output        io_cpu_s2_xcpt_ma_st,
  output        io_cpu_s2_xcpt_pf_ld,
  output        io_cpu_s2_xcpt_pf_st,
  output        io_cpu_s2_xcpt_ae_ld,
  output        io_cpu_s2_xcpt_ae_st,
  input         io_cpu_invalidate_lr,
  output        io_cpu_ordered,
  output        io_ptw_req_valid,
  output [19:0] io_ptw_req_bits_addr,
  input         io_ptw_resp_valid,
  input  [1:0]  io_ptw_status_dprv,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_mem_0_a_ready,
  output        io_mem_0_a_valid,
  output [2:0]  io_mem_0_a_bits_opcode,
  output [2:0]  io_mem_0_a_bits_param,
  output [3:0]  io_mem_0_a_bits_size,
  output [31:0] io_mem_0_a_bits_address,
  output [3:0]  io_mem_0_a_bits_mask,
  output [31:0] io_mem_0_a_bits_data,
  output        io_mem_0_b_ready,
  input         io_mem_0_b_valid,
  input  [1:0]  io_mem_0_b_bits_param,
  input  [31:0] io_mem_0_b_bits_address,
  input         io_mem_0_c_ready,
  output        io_mem_0_c_valid,
  output [31:0] io_mem_0_c_bits_address,
  output        io_mem_0_d_ready,
  input         io_mem_0_d_valid,
  input  [2:0]  io_mem_0_d_bits_opcode,
  input  [3:0]  io_mem_0_d_bits_size,
  input         io_mem_0_d_bits_source,
  input  [31:0] io_mem_0_d_bits_data,
  input         io_mem_0_e_ready,
  output        io_mem_0_e_valid
);
  wire  metaArb_io_in_0_valid;
  wire  metaArb_io_in_0_bits_write;
  wire [7:0] metaArb_io_in_0_bits_idx;
  wire  metaArb_io_in_1_valid;
  wire  metaArb_io_in_1_bits_write;
  wire [7:0] metaArb_io_in_1_bits_idx;
  wire  metaArb_io_in_2_valid;
  wire  metaArb_io_in_2_bits_write;
  wire [7:0] metaArb_io_in_2_bits_idx;
  wire  metaArb_io_in_3_ready;
  wire  metaArb_io_in_3_valid;
  wire  metaArb_io_in_3_bits_write;
  wire [7:0] metaArb_io_in_3_bits_idx;
  wire  metaArb_io_in_4_ready;
  wire  metaArb_io_in_4_valid;
  wire  metaArb_io_in_4_bits_write;
  wire [7:0] metaArb_io_in_4_bits_idx;
  wire  metaArb_io_in_5_ready;
  wire  metaArb_io_in_5_valid;
  wire  metaArb_io_in_5_bits_write;
  wire [7:0] metaArb_io_in_5_bits_idx;
  wire  metaArb_io_in_6_ready;
  wire  metaArb_io_in_6_valid;
  wire  metaArb_io_in_6_bits_write;
  wire [7:0] metaArb_io_in_6_bits_idx;
  wire  metaArb_io_in_7_ready;
  wire  metaArb_io_in_7_valid;
  wire  metaArb_io_in_7_bits_write;
  wire [7:0] metaArb_io_in_7_bits_idx;
  wire  metaArb_io_out_ready;
  wire  metaArb_io_out_valid;
  wire  metaArb_io_out_bits_write;
  wire [7:0] metaArb_io_out_bits_idx;
  wire  data_clock;
  wire  data_io_req_valid;
  wire [13:0] data_io_req_bits_addr;
  wire  data_io_req_bits_write;
  wire [31:0] data_io_req_bits_wdata;
  wire [3:0] data_io_req_bits_eccMask;
  wire [31:0] data_io_resp_0;
  wire  dataArb_io_in_0_valid;
  wire [13:0] dataArb_io_in_0_bits_addr;
  wire  dataArb_io_in_0_bits_write;
  wire [31:0] dataArb_io_in_0_bits_wdata;
  wire [3:0] dataArb_io_in_0_bits_eccMask;
  wire  dataArb_io_in_1_ready;
  wire  dataArb_io_in_1_valid;
  wire [13:0] dataArb_io_in_1_bits_addr;
  wire  dataArb_io_in_1_bits_write;
  wire [31:0] dataArb_io_in_1_bits_wdata;
  wire [3:0] dataArb_io_in_1_bits_eccMask;
  wire  dataArb_io_in_2_ready;
  wire  dataArb_io_in_2_valid;
  wire [13:0] dataArb_io_in_2_bits_addr;
  wire  dataArb_io_in_2_bits_write;
  wire [31:0] dataArb_io_in_2_bits_wdata;
  wire [3:0] dataArb_io_in_2_bits_eccMask;
  wire  dataArb_io_in_3_ready;
  wire  dataArb_io_in_3_valid;
  wire [13:0] dataArb_io_in_3_bits_addr;
  wire  dataArb_io_in_3_bits_write;
  wire [31:0] dataArb_io_in_3_bits_wdata;
  wire [3:0] dataArb_io_in_3_bits_eccMask;
  wire  dataArb_io_out_ready;
  wire  dataArb_io_out_valid;
  wire [13:0] dataArb_io_out_bits_addr;
  wire  dataArb_io_out_bits_write;
  wire [31:0] dataArb_io_out_bits_wdata;
  wire [3:0] dataArb_io_out_bits_eccMask;
  wire [31:0] _T_117;
  wire [7:0] _T_118;
  wire [7:0] _T_119;
  wire [7:0] _T_120;
  wire [7:0] _T_121;
  wire [15:0] _T_122;
  wire [15:0] _T_123;
  wire [31:0] _T_124;
  wire  _T_133;
  reg  s1_valid;
  reg [31:0] _RAND_0;
  wire  _T_136;
  reg  s1_probe;
  reg [31:0] _RAND_1;
  reg [1:0] probe_bits_param;
  reg [31:0] _RAND_2;
  reg [31:0] probe_bits_address;
  reg [31:0] _RAND_3;
  wire [1:0] _GEN_2;
  wire [31:0] _GEN_5;
  wire  _T_144;
  wire  s1_valid_masked;
  wire  _T_146;
  wire  s1_valid_not_nacked;
  reg [31:0] s1_req_addr;
  reg [31:0] _RAND_4;
  reg [6:0] s1_req_tag;
  reg [31:0] _RAND_5;
  reg [4:0] s1_req_cmd;
  reg [31:0] _RAND_6;
  reg [2:0] s1_req_typ;
  reg [31:0] _RAND_7;
  reg  s1_req_phys;
  reg [31:0] _RAND_8;
  wire  _T_148;
  wire  _T_149;
  wire [17:0] _T_150;
  wire [5:0] _T_151;
  wire [25:0] _T_152;
  wire [31:0] _T_153;
  wire [31:0] _GEN_8;
  wire [6:0] _GEN_9;
  wire [4:0] _GEN_10;
  wire [2:0] _GEN_11;
  wire  _GEN_12;
  wire  _T_155;
  wire  _T_157;
  wire  _T_158;
  wire  _T_160;
  wire  _T_161;
  wire  _T_166;
  wire  _T_167;
  wire  _T_168;
  wire  _T_169;
  wire  _T_170;
  wire  _T_171;
  wire  _T_172;
  wire  _T_178;
  wire  _T_179;
  wire  _T_180;
  wire  _T_181;
  wire  _T_182;
  wire  _T_183;
  wire  _T_184;
  wire  _T_185;
  wire  _T_186;
  wire  _T_187;
  wire  s1_read;
  wire  _T_189;
  wire  _T_191;
  wire  _T_192;
  wire  _T_195;
  wire  s1_write;
  wire  s1_readwrite;
  wire  s1_sfence;
  reg  s1_flush_valid;
  reg [31:0] _RAND_9;
  reg  cached_grant_wait;
  reg [31:0] _RAND_10;
  reg  release_ack_wait;
  reg [31:0] _RAND_11;
  reg [2:0] release_state;
  reg [31:0] _RAND_12;
  wire  _T_232;
  wire  _T_233;
  wire  inWriteback;
  wire  _T_235;
  wire  _T_237;
  wire  _T_238;
  wire  _T_241;
  reg  uncachedInFlight_0;
  reg [31:0] _RAND_13;
  reg [31:0] uncachedReqs_0_addr;
  reg [31:0] _RAND_14;
  reg [6:0] uncachedReqs_0_tag;
  reg [31:0] _RAND_15;
  reg [2:0] uncachedReqs_0_typ;
  reg [31:0] _RAND_16;
  wire  _T_246;
  wire  _T_248;
  wire  _T_249;
  wire  _T_251;
  wire  _T_252;
  wire  _T_257;
  wire  _T_258;
  wire  _T_259;
  wire  _T_260;
  wire  _T_261;
  wire  _T_262;
  wire  _T_263;
  wire  _T_269;
  wire  _T_270;
  wire  _T_271;
  wire  _T_272;
  wire  _T_273;
  wire  _T_274;
  wire  _T_275;
  wire  _T_276;
  wire  _T_277;
  wire  _T_278;
  wire  _T_279;
  wire  _T_281;
  wire  _T_283;
  wire  _T_284;
  wire  _T_287;
  wire  _T_314;
  wire  _T_321;
  wire  s0_needsRead;
  wire  _T_356;
  wire [1:0] _T_360;
  wire  _T_364;
  wire  _T_365;
  wire  _GEN_14;
  wire [7:0] _T_375;
  wire  _T_379;
  wire  _GEN_16;
  wire  tlb_clock;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [31:0] tlb_io_req_bits_vaddr;
  wire  tlb_io_req_bits_instruction;
  wire [1:0] tlb_io_req_bits_size;
  wire [4:0] tlb_io_req_bits_cmd;
  wire  tlb_io_resp_miss;
  wire [31:0] tlb_io_resp_paddr;
  wire  tlb_io_resp_pf_ld;
  wire  tlb_io_resp_pf_st;
  wire  tlb_io_resp_pf_inst;
  wire  tlb_io_resp_ae_ld;
  wire  tlb_io_resp_ae_st;
  wire  tlb_io_resp_ae_inst;
  wire  tlb_io_resp_ma_ld;
  wire  tlb_io_resp_ma_st;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_valid;
  wire [19:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_resp_valid;
  wire [1:0] tlb_io_ptw_status_dprv;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_sum;
  wire  tlb_io_ptw_pmp_0_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a;
  wire  tlb_io_ptw_pmp_0_cfg_x;
  wire  tlb_io_ptw_pmp_0_cfg_w;
  wire  tlb_io_ptw_pmp_0_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_0_addr;
  wire [31:0] tlb_io_ptw_pmp_0_mask;
  wire  tlb_io_ptw_pmp_1_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a;
  wire  tlb_io_ptw_pmp_1_cfg_x;
  wire  tlb_io_ptw_pmp_1_cfg_w;
  wire  tlb_io_ptw_pmp_1_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_1_addr;
  wire [31:0] tlb_io_ptw_pmp_1_mask;
  wire  tlb_io_ptw_pmp_2_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a;
  wire  tlb_io_ptw_pmp_2_cfg_x;
  wire  tlb_io_ptw_pmp_2_cfg_w;
  wire  tlb_io_ptw_pmp_2_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_2_addr;
  wire [31:0] tlb_io_ptw_pmp_2_mask;
  wire  tlb_io_ptw_pmp_3_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a;
  wire  tlb_io_ptw_pmp_3_cfg_x;
  wire  tlb_io_ptw_pmp_3_cfg_w;
  wire  tlb_io_ptw_pmp_3_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_3_addr;
  wire [31:0] tlb_io_ptw_pmp_3_mask;
  wire  tlb_io_ptw_pmp_4_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a;
  wire  tlb_io_ptw_pmp_4_cfg_x;
  wire  tlb_io_ptw_pmp_4_cfg_w;
  wire  tlb_io_ptw_pmp_4_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_4_addr;
  wire [31:0] tlb_io_ptw_pmp_4_mask;
  wire  tlb_io_ptw_pmp_5_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a;
  wire  tlb_io_ptw_pmp_5_cfg_x;
  wire  tlb_io_ptw_pmp_5_cfg_w;
  wire  tlb_io_ptw_pmp_5_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_5_addr;
  wire [31:0] tlb_io_ptw_pmp_5_mask;
  wire  tlb_io_ptw_pmp_6_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a;
  wire  tlb_io_ptw_pmp_6_cfg_x;
  wire  tlb_io_ptw_pmp_6_cfg_w;
  wire  tlb_io_ptw_pmp_6_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_6_addr;
  wire [31:0] tlb_io_ptw_pmp_6_mask;
  wire  tlb_io_ptw_pmp_7_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a;
  wire  tlb_io_ptw_pmp_7_cfg_x;
  wire  tlb_io_ptw_pmp_7_cfg_w;
  wire  tlb_io_ptw_pmp_7_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_7_addr;
  wire [31:0] tlb_io_ptw_pmp_7_mask;
  wire  _T_384;
  wire  _T_385;
  wire  _T_390;
  wire  _T_392;
  wire  _T_393;
  wire  _T_395;
  wire  _T_396;
  wire  _GEN_17;
  wire  _T_398;
  wire  _T_399;
  wire  _T_408;
  wire [32:0] _T_410;
  wire [31:0] _T_411;
  wire  _T_412;
  wire  s1_hit_way;
  wire [1:0] s1_hit_state_state;
  wire [1:0] _T_428;
  wire  _T_430;
  wire  _T_434;
  wire  _T_438;
  wire  _T_441;
  wire [1:0] _T_442;
  wire  _T_443;
  wire [1:0] _T_445;
  wire  _T_447;
  wire [1:0] _T_450;
  wire [1:0] _T_451;
  wire [1:0] _T_454;
  wire [3:0] _T_455;
  wire [3:0] s1_mask;
  wire  _T_457;
  wire  _T_458;
  reg  _T_461;
  reg [31:0] _RAND_17;
  wire [1:0] _T_462;
  wire [2:0] _T_463;
  wire [1:0] _T_464;
  wire [2:0] _T_465;
  wire [5:0] _T_466;
  wire  _T_468;
  wire  _T_470;
  wire  s2_valid;
  reg  s2_probe;
  reg [31:0] _RAND_18;
  wire  _T_473;
  wire  _T_474;
  wire  releaseInFlight;
  reg  _T_478;
  reg [31:0] _RAND_19;
  wire  s2_valid_masked;
  reg [31:0] s2_req_addr;
  reg [31:0] _RAND_20;
  reg [6:0] s2_req_tag;
  reg [31:0] _RAND_21;
  reg [4:0] s2_req_cmd;
  reg [31:0] _RAND_22;
  reg [2:0] s2_req_typ;
  reg [31:0] _RAND_23;
  reg  s2_req_phys;
  reg [31:0] _RAND_24;
  wire [25:0] _T_479;
  wire [31:0] _GEN_234;
  wire [31:0] acquire_address;
  reg  s2_uncached;
  reg [31:0] _RAND_25;
  wire  _T_482;
  wire [31:0] _GEN_19;
  wire [6:0] _GEN_20;
  wire [4:0] _GEN_21;
  wire [2:0] _GEN_22;
  wire  _GEN_23;
  wire  _GEN_25;
  wire  _T_488;
  wire  _T_490;
  wire  _T_491;
  wire  _T_493;
  wire  _T_494;
  wire  _T_499;
  wire  _T_500;
  wire  _T_501;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_511;
  wire  _T_512;
  wire  _T_513;
  wire  _T_514;
  wire  _T_515;
  wire  _T_516;
  wire  _T_517;
  wire  _T_518;
  wire  _T_519;
  wire  _T_520;
  wire  s2_read;
  wire  _T_522;
  wire  _T_524;
  wire  _T_525;
  wire  _T_528;
  wire  s2_write;
  wire  s2_readwrite;
  reg  s2_flush_valid_pre_tag_ecc;
  reg [31:0] _RAND_26;
  wire  _T_571;
  reg [31:0] s2_data;
  reg [31:0] _RAND_27;
  wire [31:0] _GEN_27;
  reg [1:0] s2_probe_state_state;
  reg [31:0] _RAND_28;
  wire [1:0] _GEN_29;
  reg [1:0] s2_hit_state_state;
  reg [31:0] _RAND_29;
  wire [1:0] _GEN_31;
  reg  s2_waw_hazard;
  reg [31:0] _RAND_30;
  wire  _GEN_32;
  wire  s2_hit_valid;
  wire  _T_651;
  wire  _T_652;
  wire  _T_655;
  wire [1:0] _T_656;
  wire [3:0] _T_657;
  wire  _T_744;
  wire [1:0] _T_746;
  wire  _T_747;
  wire [1:0] _T_749;
  wire  _T_750;
  wire [1:0] _T_752;
  wire  _T_753;
  wire [1:0] _T_755;
  wire  _T_756;
  wire [1:0] _T_758;
  wire  _T_759;
  wire [1:0] _T_761;
  wire  _T_762;
  wire  _T_763;
  wire [1:0] _T_764;
  wire  _T_765;
  wire  _T_766;
  wire [1:0] _T_767;
  wire  _T_768;
  wire  _T_769;
  wire [1:0] _T_770;
  wire  _T_771;
  wire  _T_772;
  wire [1:0] _T_773;
  wire  _T_774;
  wire  _T_775;
  wire [1:0] _T_776;
  wire  _T_777;
  wire  s2_hit;
  wire [1:0] s2_grow_param;
  wire [7:0] _T_779;
  wire [7:0] _T_780;
  wire [7:0] _T_781;
  wire [7:0] _T_782;
  wire [1:0] _T_855;
  wire [15:0] _T_876;
  wire [15:0] _T_877;
  wire [31:0] s2_data_corrected;
  wire  _T_880;
  wire  s2_valid_hit_pre_data_ecc;
  wire  _T_888;
  wire  s2_valid_hit;
  wire  _T_895;
  wire  _T_896;
  wire  _T_898;
  wire  s2_valid_miss;
  wire  _T_900;
  wire  _T_901;
  wire  _T_905;
  wire  s2_valid_cached_miss;
  wire  s2_valid_uncached;
  wire  _T_910;
  wire  _T_911;
  reg [1:0] _T_926_state;
  reg [31:0] _RAND_31;
  wire [1:0] _GEN_35;
  wire [1:0] s2_victim_state_state;
  wire [3:0] _T_927;
  wire  _T_1015;
  wire  _T_1019;
  wire  _T_1020;
  wire  _T_1023;
  wire  _T_1024;
  wire  _T_1027;
  wire  _T_1028;
  wire  _T_1031;
  wire  _T_1032;
  wire  _T_1035;
  wire  _T_1036;
  wire  _T_1039;
  wire  _T_1040;
  wire  _T_1043;
  wire  _T_1044;
  wire  _T_1047;
  wire  s2_prb_ack_data;
  wire [3:0] _T_1064;
  wire  _T_1152;
  wire  _T_1156;
  wire  _T_1157;
  wire  _T_1160;
  wire  _T_1161;
  wire  _T_1164;
  wire  _T_1165;
  wire  _T_1168;
  wire  _T_1169;
  wire  _T_1172;
  wire  _T_1173;
  wire  _T_1176;
  wire  _T_1177;
  wire  _T_1180;
  wire  _T_1181;
  wire  _T_1184;
  wire  s2_victim_dirty;
  wire  _T_1187;
  wire  s2_update_meta;
  wire  _T_1190;
  wire  _T_1191;
  wire  _T_1192;
  wire  _T_1193;
  wire  _T_1195;
  wire  _T_1197;
  wire  _T_1198;
  wire  _T_1200;
  wire  _T_1201;
  wire  _T_1202;
  wire  _T_1203;
  wire  _GEN_36;
  wire [31:0] _T_1214;
  wire [7:0] _T_1215;
  wire  _T_1219;
  wire [7:0] _T_1223;
  reg [4:0] lrscCount;
  reg [31:0] _RAND_32;
  wire  lrscValid;
  wire  _T_1248;
  wire [5:0] _T_1250;
  wire [5:0] _T_1251;
  wire [4:0] _T_1252;
  wire [4:0] _GEN_39;
  wire  _T_1255;
  wire  _T_1256;
  wire [4:0] _GEN_40;
  wire  _T_1262;
  reg [4:0] pstore1_cmd;
  reg [31:0] _RAND_33;
  wire [4:0] _GEN_41;
  reg [31:0] pstore1_addr;
  reg [31:0] _RAND_34;
  wire [31:0] _GEN_42;
  reg [31:0] a_data;
  reg [31:0] _RAND_35;
  wire [31:0] _GEN_43;
  reg [3:0] pstore1_mask;
  reg [31:0] _RAND_36;
  wire [3:0] _GEN_45;
  wire  _T_1350;
  wire  _T_1351;
  reg  _T_1354;
  reg [31:0] _RAND_37;
  wire  _GEN_46;
  reg  pstore2_valid;
  reg [31:0] _RAND_38;
  wire  _T_1358;
  wire  _T_1359;
  wire  _T_1360;
  wire  pstore_drain_structural;
  wire  pstore_drain_opportunistic;
  wire  pstore_drain_on_miss;
  wire  _T_1368;
  wire  _T_1369;
  wire  _T_1370;
  wire  _T_1371;
  wire  _T_1372;
  wire  _T_1373;
  wire  _T_1374;
  reg  _T_1379;
  reg [31:0] _RAND_39;
  wire  _T_1381;
  wire  _T_1383;
  wire  _T_1384;
  wire  _T_1385;
  wire  _T_1387;
  wire  _T_1391;
  wire  _T_1392;
  wire  _T_1394;
  wire  _T_1395;
  wire  _T_1396;
  wire  _T_1398;
  wire  advance_pstore1;
  wire  _T_1401;
  wire  _T_1402;
  reg [31:0] pstore2_addr;
  reg [31:0] _RAND_40;
  wire [31:0] _GEN_47;
  wire [11:0] _T_1408;
  wire [7:0] _T_1417;
  wire  _T_1418;
  reg [7:0] _T_1422;
  reg [31:0] _RAND_41;
  wire [7:0] _GEN_49;
  wire [7:0] _T_1423;
  wire  _T_1424;
  reg [7:0] _T_1428;
  reg [31:0] _RAND_42;
  wire [7:0] _GEN_50;
  wire [7:0] _T_1429;
  wire  _T_1430;
  reg [7:0] _T_1434;
  reg [31:0] _RAND_43;
  wire [7:0] _GEN_51;
  wire [7:0] _T_1435;
  wire  _T_1436;
  reg [7:0] _T_1440;
  reg [31:0] _RAND_44;
  wire [7:0] _GEN_52;
  wire [15:0] _T_1441;
  wire [15:0] _T_1442;
  wire [31:0] pstore2_storegen_data;
  reg [3:0] pstore2_storegen_mask;
  reg [31:0] _RAND_45;
  wire [3:0] _T_1449;
  wire [3:0] _T_1451;
  wire [3:0] _GEN_53;
  wire [31:0] _T_1453;
  wire [31:0] _T_1455;
  wire [3:0] _T_1460;
  wire  _T_1461;
  wire  _T_1462;
  wire  _T_1463;
  wire  _T_1464;
  wire [1:0] _T_1473;
  wire [1:0] _T_1474;
  wire [3:0] _T_1475;
  wire [11:0] _T_1476;
  wire [11:0] _T_1477;
  wire  _T_1478;
  wire [1:0] _T_1491;
  wire [1:0] _T_1492;
  wire [3:0] _T_1493;
  wire  _T_1494;
  wire  _T_1495;
  wire  _T_1496;
  wire  _T_1497;
  wire [1:0] _T_1498;
  wire [1:0] _T_1499;
  wire [3:0] _T_1500;
  wire  _T_1501;
  wire  _T_1502;
  wire  _T_1503;
  wire  _T_1504;
  wire [1:0] _T_1513;
  wire [1:0] _T_1514;
  wire [3:0] _T_1515;
  wire  _T_1516;
  wire  _T_1517;
  wire  _T_1518;
  wire  _T_1519;
  wire [1:0] _T_1520;
  wire [1:0] _T_1521;
  wire [3:0] _T_1522;
  wire [3:0] _T_1523;
  wire  _T_1525;
  wire [3:0] _T_1526;
  wire  _T_1528;
  wire  _T_1529;
  wire  _T_1530;
  wire  _T_1531;
  wire  _T_1534;
  wire  _T_1535;
  wire  _T_1536;
  wire  _T_1537;
  wire  _T_1538;
  wire [1:0] _T_1547;
  wire [1:0] _T_1548;
  wire [3:0] _T_1549;
  wire  _T_1550;
  wire  _T_1551;
  wire  _T_1552;
  wire  _T_1553;
  wire [1:0] _T_1554;
  wire [1:0] _T_1555;
  wire [3:0] _T_1556;
  wire [3:0] _T_1579;
  wire  _T_1581;
  wire [3:0] _T_1582;
  wire  _T_1584;
  wire  _T_1585;
  wire  _T_1586;
  wire  _T_1587;
  wire  s1_hazard;
  wire  s1_raw_hazard;
  wire  _T_1592;
  wire  _GEN_54;
  wire [2:0] acquire__param;
  wire [3:0] get_size;
  wire  _T_1799;
  wire [1:0] _T_1801;
  wire [1:0] _T_1804;
  wire  _T_1806;
  wire  _T_1808;
  wire  _T_1809;
  wire  _T_1811;
  wire  _T_1813;
  wire  _T_1814;
  wire  _T_1816;
  wire  _T_1817;
  wire  _T_1818;
  wire  _T_1819;
  wire  _T_1821;
  wire  _T_1822;
  wire  _T_1823;
  wire  _T_1824;
  wire  _T_1825;
  wire  _T_1826;
  wire  _T_1827;
  wire  _T_1828;
  wire  _T_1829;
  wire  _T_1830;
  wire  _T_1831;
  wire  _T_1832;
  wire  _T_1833;
  wire [1:0] _T_1834;
  wire [1:0] _T_1835;
  wire [3:0] _T_1836;
  wire [3:0] put_size;
  wire [3:0] _T_2060_size;
  wire [3:0] _T_2187_size;
  wire [3:0] _T_2314_size;
  wire [3:0] _T_2441_size;
  wire [3:0] _T_2568_size;
  wire [3:0] _T_2695_size;
  wire [3:0] _T_2822_size;
  wire [3:0] _T_2949_size;
  wire [3:0] _T_3076_size;
  wire  _T_3116;
  wire [2:0] _T_3117_opcode;
  wire [2:0] _T_3117_param;
  wire [3:0] _T_3117_size;
  wire [31:0] _T_3117_address;
  wire [3:0] _T_3117_mask;
  wire [31:0] _T_3117_data;
  wire  _T_3118;
  wire [2:0] _T_3119_opcode;
  wire [2:0] _T_3119_param;
  wire [3:0] _T_3119_size;
  wire [31:0] _T_3119_address;
  wire [3:0] _T_3119_mask;
  wire [31:0] _T_3119_data;
  wire  _T_3120;
  wire [2:0] _T_3121_opcode;
  wire [2:0] _T_3121_param;
  wire [3:0] _T_3121_size;
  wire [31:0] _T_3121_address;
  wire [3:0] _T_3121_mask;
  wire [31:0] _T_3121_data;
  wire  _T_3122;
  wire [2:0] _T_3123_opcode;
  wire [2:0] _T_3123_param;
  wire [3:0] _T_3123_size;
  wire [31:0] _T_3123_address;
  wire [3:0] _T_3123_mask;
  wire [31:0] _T_3123_data;
  wire  _T_3124;
  wire [2:0] _T_3125_opcode;
  wire [2:0] _T_3125_param;
  wire [3:0] _T_3125_size;
  wire [31:0] _T_3125_address;
  wire [3:0] _T_3125_mask;
  wire [31:0] _T_3125_data;
  wire  _T_3126;
  wire [2:0] _T_3127_opcode;
  wire [2:0] _T_3127_param;
  wire [3:0] _T_3127_size;
  wire [31:0] _T_3127_address;
  wire [3:0] _T_3127_mask;
  wire [31:0] _T_3127_data;
  wire  _T_3128;
  wire [2:0] _T_3129_opcode;
  wire [2:0] _T_3129_param;
  wire [3:0] _T_3129_size;
  wire [31:0] _T_3129_address;
  wire [3:0] _T_3129_mask;
  wire [31:0] _T_3129_data;
  wire  _T_3130;
  wire [2:0] _T_3131_opcode;
  wire [2:0] _T_3131_param;
  wire [3:0] _T_3131_size;
  wire [31:0] _T_3131_address;
  wire [3:0] _T_3131_mask;
  wire [31:0] _T_3131_data;
  wire  _T_3132;
  wire [2:0] atomics_opcode;
  wire [2:0] atomics_param;
  wire [3:0] atomics_size;
  wire [31:0] atomics_address;
  wire [3:0] atomics_mask;
  wire [31:0] atomics_data;
  wire  _T_3137;
  wire  _T_3143;
  wire  _T_3144;
  wire  _T_3148;
  wire  _T_3150;
  wire [2:0] _T_3151_opcode;
  wire [2:0] _T_3151_param;
  wire [3:0] _T_3151_size;
  wire [31:0] _T_3151_address;
  wire [3:0] _T_3151_mask;
  wire [31:0] _T_3151_data;
  wire [2:0] _T_3152_opcode;
  wire [2:0] _T_3152_param;
  wire [3:0] _T_3152_size;
  wire [31:0] _T_3152_address;
  wire [3:0] _T_3152_mask;
  wire [31:0] _T_3152_data;
  wire [2:0] _T_3153_opcode;
  wire [2:0] _T_3153_param;
  wire [3:0] _T_3153_size;
  wire [31:0] _T_3153_address;
  wire [3:0] _T_3153_mask;
  wire [31:0] _T_3153_data;
  wire  _T_3157;
  wire  _T_3158;
  wire  _GEN_55;
  wire [31:0] _GEN_56;
  wire [6:0] _GEN_57;
  wire [2:0] _GEN_59;
  wire  _GEN_62;
  wire [31:0] _GEN_63;
  wire [6:0] _GEN_64;
  wire [2:0] _GEN_66;
  wire  _GEN_69;
  wire  _GEN_70;
  wire [31:0] _GEN_71;
  wire [6:0] _GEN_72;
  wire [2:0] _GEN_74;
  wire  _GEN_77;
  wire  _T_3164;
  wire [26:0] _T_3167;
  wire [11:0] _T_3168;
  wire [11:0] _T_3169;
  wire [9:0] _T_3170;
  wire  _T_3171;
  wire [9:0] _T_3173;
  reg [9:0] _T_3176;
  reg [31:0] _RAND_46;
  wire [10:0] _T_3178;
  wire [10:0] _T_3179;
  wire [9:0] _T_3180;
  wire  d_first;
  wire  _T_3183;
  wire  _T_3185;
  wire  d_last;
  wire  d_done;
  wire [9:0] _T_3186;
  wire [9:0] _T_3187;
  wire [9:0] _T_3188;
  wire [9:0] _GEN_78;
  wire [11:0] _GEN_235;
  wire [11:0] d_address_inc;
  wire  _T_3191;
  wire  _T_3192;
  wire  grantIsCached;
  wire  _T_3196;
  wire  _T_3197;
  wire  _T_3198;
  wire  _T_3199;
  wire  grantIsUncached;
  wire  grantIsVoluntary;
  reg  grantInProgress;
  reg [31:0] _RAND_47;
  reg [2:0] blockProbeAfterGrantCount;
  reg [31:0] _RAND_48;
  wire  _T_3208;
  wire [3:0] _T_3210;
  wire [3:0] _T_3211;
  wire [2:0] _T_3212;
  wire [2:0] _GEN_79;
  wire  _T_3214;
  wire  _T_3215;
  wire  _T_3218;
  wire  _T_3221;
  wire  _T_3223;
  wire  _GEN_80;
  wire  _GEN_81;
  wire [2:0] _GEN_82;
  wire  _GEN_84;
  wire  _GEN_85;
  wire [2:0] _GEN_86;
  wire  _T_3229;
  wire  _T_3230;
  wire [1:0] _T_3233;
  wire  _T_3234;
  wire  _T_3238;
  wire  _T_3239;
  wire  _T_3241;
  wire  _GEN_88;
  wire [7:0] _T_3243;
  wire [7:0] _T_3244;
  wire [7:0] _T_3245;
  wire [7:0] _T_3246;
  wire [15:0] _T_3247;
  wire [15:0] _T_3248;
  wire [31:0] _T_3249;
  wire [29:0] _T_3251;
  wire [1:0] _T_3252;
  wire [31:0] _T_3253;
  wire [31:0] _GEN_89;
  wire [4:0] _GEN_90;
  wire [2:0] _GEN_91;
  wire [6:0] _GEN_92;
  wire [31:0] _GEN_93;
  wire  _GEN_95;
  wire [31:0] _GEN_96;
  wire [4:0] _GEN_97;
  wire [2:0] _GEN_98;
  wire [6:0] _GEN_99;
  wire [31:0] _GEN_100;
  wire  _T_3257;
  wire  _T_3258;
  wire  _T_3259;
  wire  _T_3260;
  wire  _T_3262;
  wire  _GEN_102;
  wire  _GEN_103;
  wire  _GEN_104;
  wire [2:0] _GEN_105;
  wire  _GEN_107;
  wire [31:0] _GEN_108;
  wire [4:0] _GEN_109;
  wire [2:0] _GEN_110;
  wire [6:0] _GEN_111;
  wire [31:0] _GEN_112;
  wire  _GEN_114;
  wire  _T_3264;
  wire  _T_3267;
  wire  _T_3268;
  wire  _GEN_115;
  wire [31:0] _GEN_236;
  wire [31:0] _T_3271;
  wire  _T_3276;
  wire  _T_3278;
  wire  _T_3279;
  wire  _T_3280;
  wire  _T_3282;
  reg  blockUncachedGrant;
  reg [31:0] _RAND_49;
  wire  _T_3400;
  wire  _T_3401;
  wire  _GEN_116;
  wire  _GEN_117;
  wire  _GEN_118;
  wire  _GEN_119;
  wire  _GEN_120;
  wire  _GEN_121;
  wire  _GEN_122;
  wire  _GEN_123;
  wire  _GEN_124;
  wire  _T_3408;
  wire  _T_3409;
  wire  _T_3413;
  wire  _T_3415;
  wire  _T_3417;
  wire  _T_3418;
  wire  _T_3421;
  wire  _T_3422;
  wire  _T_3425;
  wire  _T_3426;
  wire  _T_3429;
  wire  _T_3431;
  wire  _T_3432;
  wire  _T_3434;
  wire  _T_3435;
  wire  _T_3436;
  wire [7:0] _T_3438;
  wire  _T_3441;
  reg [9:0] _T_3454;
  reg [31:0] _RAND_50;
  wire [10:0] _T_3456;
  wire [10:0] _T_3457;
  wire [9:0] _T_3458;
  wire  c_first;
  wire [9:0] _T_3465;
  wire [9:0] _GEN_125;
  wire  _T_3467;
  wire  releaseRejected;
  wire  _T_3468;
  reg  s1_release_data_valid;
  reg [31:0] _RAND_51;
  wire  _T_3471;
  wire  _T_3472;
  reg  s2_release_data_valid;
  reg [31:0] _RAND_52;
  wire [1:0] _T_3478;
  wire [1:0] _GEN_237;
  wire [2:0] _T_3479;
  wire [1:0] _T_3480;
  wire [1:0] _T_3481;
  wire [10:0] _GEN_238;
  wire [11:0] _T_3482;
  wire [10:0] releaseDataBeat;
  wire [2:0] _GEN_129;
  wire  _T_3517;
  wire  _T_3521;
  wire  _T_3523;
  wire [2:0] _T_3525;
  wire  _GEN_130;
  wire [2:0] _GEN_138;
  wire  _T_3532;
  wire  _T_3533;
  wire  _T_3536;
  wire [2:0] _T_3537;
  wire  _GEN_139;
  wire  _GEN_140;
  wire [2:0] _GEN_141;
  wire  _GEN_142;
  wire [2:0] _GEN_143;
  wire  _GEN_144;
  wire  _GEN_152;
  wire  _T_3539;
  wire [7:0] _T_3541;
  wire [2:0] _GEN_153;
  wire  _GEN_154;
  wire  _GEN_155;
  wire [7:0] _GEN_156;
  wire [2:0] _GEN_157;
  wire  _GEN_158;
  wire  _T_3543;
  wire [2:0] _GEN_159;
  wire  _GEN_160;
  wire [2:0] _GEN_161;
  wire  _T_3545;
  wire [2:0] _GEN_162;
  wire  _GEN_163;
  wire [2:0] _GEN_171;
  wire [2:0] _GEN_172;
  wire [2:0] _GEN_180;
  wire  _T_3549;
  wire  _T_3550;
  wire [2:0] _GEN_181;
  wire  _T_3636;
  wire  _GEN_182;
  wire [2:0] _GEN_192;
  wire  _GEN_193;
  wire  _T_3639;
  wire  _T_3640;
  wire [3:0] _T_3642;
  wire [5:0] _GEN_246;
  wire [5:0] _T_3643;
  wire [31:0] _GEN_247;
  wire [31:0] _T_3644;
  wire  _T_3650;
  wire  _T_3651;
  wire [7:0] _T_3653;
  wire  _T_3655;
  wire [2:0] _GEN_194;
  wire  _T_3657;
  wire  _T_3658;
  wire  _T_3661;
  wire  _T_3663;
  wire  s1_xcpt_valid;
  reg  _T_3667;
  reg [31:0] _RAND_53;
  reg  _T_3669_pf_ld;
  reg [31:0] _RAND_54;
  reg  _T_3669_pf_st;
  reg [31:0] _RAND_55;
  reg  _T_3669_ae_ld;
  reg [31:0] _RAND_56;
  reg  _T_3669_ae_st;
  reg [31:0] _RAND_57;
  reg  _T_3669_ma_ld;
  reg [31:0] _RAND_58;
  reg  _T_3669_ma_st;
  reg [31:0] _RAND_59;
  wire  _GEN_197;
  wire  _GEN_198;
  wire  _GEN_200;
  wire  _GEN_201;
  wire  _GEN_203;
  wire  _GEN_204;
  wire  _T_3687_pf_ld;
  wire  _T_3687_pf_st;
  wire  _T_3687_ae_ld;
  wire  _T_3687_ae_st;
  wire  _T_3687_ma_ld;
  wire  _T_3687_ma_st;
  wire  _T_3690;
  wire  _T_3691;
  wire  _T_3693;
  wire  _GEN_207;
  wire  _GEN_208;
  wire  _GEN_209;
  wire  _GEN_210;
  wire  _GEN_211;
  wire  _GEN_212;
  wire  _T_3709;
  wire  _T_3710;
  wire  _T_3712;
  wire  _T_3713;
  wire  _T_3715;
  wire  _T_3717;
  reg  doUncachedResp;
  reg [31:0] _RAND_60;
  wire  _T_3721;
  wire  _T_3723;
  wire  _GEN_213;
  wire  _T_3726;
  wire  _T_3728;
  wire [15:0] _T_3731;
  wire [15:0] _T_3732;
  wire [15:0] _T_3733;
  wire  _T_3739;
  wire  _T_3741;
  wire  _T_3742;
  wire [15:0] _T_3746;
  wire [15:0] _T_3748;
  wire [31:0] _T_3749;
  wire [7:0] _T_3751;
  wire [7:0] _T_3752;
  wire [7:0] _T_3753;
  wire  _T_3759;
  wire  _T_3761;
  wire  _T_3762;
  wire [23:0] _T_3766;
  wire [23:0] _T_3767;
  wire [23:0] _T_3768;
  wire [31:0] _T_3769;
  wire [3:0] AMOALU_io_mask;
  wire [4:0] AMOALU_io_cmd;
  wire [31:0] AMOALU_io_lhs;
  wire [31:0] AMOALU_io_rhs;
  wire [31:0] AMOALU_io_out;
  wire [31:0] _GEN_216;
  reg  resetting;
  reg [31:0] _RAND_61;
  reg  flushed;
  reg [31:0] _RAND_62;
  reg  flushing;
  reg [31:0] _RAND_63;
  reg [7:0] flushCounter;
  reg [31:0] _RAND_64;
  wire [8:0] flushCounterNext;
  wire  _T_3780;
  wire  _T_3785;
  wire  _GEN_217;
  wire  _T_3788;
  wire  _T_3789;
  wire  _T_3791;
  wire  _T_3800;
  wire  _GEN_218;
  wire  _GEN_219;
  wire  _GEN_220;
  wire  _T_3801;
  wire  _T_3803;
  wire  _T_3804;
  wire  _T_3807;
  wire  _T_3809;
  wire  _T_3812;
  wire  _GEN_221;
  wire [8:0] _GEN_222;
  wire  _GEN_223;
  wire  _T_3819;
  wire  _T_3822;
  wire  _GEN_224;
  wire [8:0] _GEN_226;
  wire  _GEN_227;
  wire  _GEN_228;
  wire  _GEN_229;
  wire [8:0] _GEN_230;
  wire  _GEN_231;
  wire  _GEN_248;
  wire  _GEN_250;
  wire  _GEN_251;
  wire  _GEN_254;
  Arbiter metaArb (
    .io_in_0_valid(metaArb_io_in_0_valid),
    .io_in_0_bits_write(metaArb_io_in_0_bits_write),
    .io_in_0_bits_idx(metaArb_io_in_0_bits_idx),
    .io_in_1_valid(metaArb_io_in_1_valid),
    .io_in_1_bits_write(metaArb_io_in_1_bits_write),
    .io_in_1_bits_idx(metaArb_io_in_1_bits_idx),
    .io_in_2_valid(metaArb_io_in_2_valid),
    .io_in_2_bits_write(metaArb_io_in_2_bits_write),
    .io_in_2_bits_idx(metaArb_io_in_2_bits_idx),
    .io_in_3_ready(metaArb_io_in_3_ready),
    .io_in_3_valid(metaArb_io_in_3_valid),
    .io_in_3_bits_write(metaArb_io_in_3_bits_write),
    .io_in_3_bits_idx(metaArb_io_in_3_bits_idx),
    .io_in_4_ready(metaArb_io_in_4_ready),
    .io_in_4_valid(metaArb_io_in_4_valid),
    .io_in_4_bits_write(metaArb_io_in_4_bits_write),
    .io_in_4_bits_idx(metaArb_io_in_4_bits_idx),
    .io_in_5_ready(metaArb_io_in_5_ready),
    .io_in_5_valid(metaArb_io_in_5_valid),
    .io_in_5_bits_write(metaArb_io_in_5_bits_write),
    .io_in_5_bits_idx(metaArb_io_in_5_bits_idx),
    .io_in_6_ready(metaArb_io_in_6_ready),
    .io_in_6_valid(metaArb_io_in_6_valid),
    .io_in_6_bits_write(metaArb_io_in_6_bits_write),
    .io_in_6_bits_idx(metaArb_io_in_6_bits_idx),
    .io_in_7_ready(metaArb_io_in_7_ready),
    .io_in_7_valid(metaArb_io_in_7_valid),
    .io_in_7_bits_write(metaArb_io_in_7_bits_write),
    .io_in_7_bits_idx(metaArb_io_in_7_bits_idx),
    .io_out_ready(metaArb_io_out_ready),
    .io_out_valid(metaArb_io_out_valid),
    .io_out_bits_write(metaArb_io_out_bits_write),
    .io_out_bits_idx(metaArb_io_out_bits_idx)
  );
  DCacheDataArray data (
    .clock(data_clock),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_eccMask(data_io_req_bits_eccMask),
    .io_resp_0(data_io_resp_0)
  );
  Arbiter_1 dataArb (
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_eccMask(dataArb_io_in_0_bits_eccMask),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_1_bits_eccMask(dataArb_io_in_1_bits_eccMask),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_write(dataArb_io_in_2_bits_write),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_2_bits_eccMask(dataArb_io_in_2_bits_eccMask),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_write(dataArb_io_in_3_bits_write),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_eccMask(dataArb_io_in_3_bits_eccMask),
    .io_out_ready(dataArb_io_out_ready),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_eccMask(dataArb_io_out_bits_eccMask)
  );
  TLB tlb (
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_size(tlb_io_req_bits_size),
    .io_req_bits_cmd(tlb_io_req_bits_cmd),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_ld(tlb_io_resp_pf_ld),
    .io_resp_pf_st(tlb_io_resp_pf_st),
    .io_resp_pf_inst(tlb_io_resp_pf_inst),
    .io_resp_ae_ld(tlb_io_resp_ae_ld),
    .io_resp_ae_st(tlb_io_resp_ae_st),
    .io_resp_ae_inst(tlb_io_resp_ae_inst),
    .io_resp_ma_ld(tlb_io_resp_ma_ld),
    .io_resp_ma_st(tlb_io_resp_ma_st),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_status_dprv(tlb_io_ptw_status_dprv),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_sum(tlb_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask)
  );
  AMOALU AMOALU (
    .io_mask(AMOALU_io_mask),
    .io_cmd(AMOALU_io_cmd),
    .io_lhs(AMOALU_io_lhs),
    .io_rhs(AMOALU_io_rhs),
    .io_out(AMOALU_io_out)
  );
  assign io_cpu_req_ready = _GEN_121;
  assign io_cpu_s2_nack = _GEN_219;
  assign io_cpu_resp_valid = _GEN_213;
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_data = _T_3769;
  assign io_cpu_resp_bits_replay = doUncachedResp;
  assign io_cpu_resp_bits_has_data = s2_read;
  assign io_cpu_resp_bits_data_word_bypass = s2_data_corrected;
  assign io_cpu_resp_bits_data_raw = s2_data_corrected;
  assign io_cpu_replay_next = _T_3717;
  assign io_cpu_s2_xcpt_ma_ld = _GEN_207;
  assign io_cpu_s2_xcpt_ma_st = _GEN_208;
  assign io_cpu_s2_xcpt_pf_ld = _GEN_209;
  assign io_cpu_s2_xcpt_pf_st = _GEN_210;
  assign io_cpu_s2_xcpt_ae_ld = _GEN_211;
  assign io_cpu_s2_xcpt_ae_st = _GEN_212;
  assign io_cpu_ordered = _T_3663;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_mem_0_a_valid = _T_3144;
  assign io_mem_0_a_bits_opcode = _T_3153_opcode;
  assign io_mem_0_a_bits_param = _T_3153_param;
  assign io_mem_0_a_bits_size = _T_3153_size;
  assign io_mem_0_a_bits_address = _T_3153_address;
  assign io_mem_0_a_bits_mask = _T_3153_mask;
  assign io_mem_0_a_bits_data = _T_3153_data;
  assign io_mem_0_b_ready = _T_3436;
  assign io_mem_0_c_valid = _GEN_163;
  assign io_mem_0_c_bits_address = probe_bits_address;
  assign io_mem_0_d_ready = _GEN_120;
  assign io_mem_0_e_valid = _T_3409;
  assign metaArb_io_in_0_valid = resetting;
  assign metaArb_io_in_0_bits_write = 1'h1;
  assign metaArb_io_in_0_bits_idx = flushCounter;
  assign metaArb_io_in_1_valid = 1'h0;
  assign metaArb_io_in_1_bits_write = 1'h1;
  assign metaArb_io_in_1_bits_idx = _T_1215;
  assign metaArb_io_in_2_valid = _T_1202;
  assign metaArb_io_in_2_bits_write = 1'h1;
  assign metaArb_io_in_2_bits_idx = _T_1223;
  assign metaArb_io_in_3_valid = _T_3276;
  assign metaArb_io_in_3_bits_write = 1'h1;
  assign metaArb_io_in_3_bits_idx = _T_1223;
  assign metaArb_io_in_4_valid = _T_3651;
  assign metaArb_io_in_4_bits_write = 1'h1;
  assign metaArb_io_in_4_bits_idx = _T_3653;
  assign metaArb_io_in_5_valid = flushing;
  assign metaArb_io_in_5_bits_write = 1'h0;
  assign metaArb_io_in_5_bits_idx = flushCounter;
  assign metaArb_io_in_6_valid = _GEN_155;
  assign metaArb_io_in_6_bits_write = 1'h0;
  assign metaArb_io_in_6_bits_idx = _GEN_156;
  assign metaArb_io_in_7_valid = io_cpu_req_valid;
  assign metaArb_io_in_7_bits_write = 1'h0;
  assign metaArb_io_in_7_bits_idx = _T_375;
  assign metaArb_io_out_ready = 1'h1;
  assign data_clock = clock;
  assign data_io_req_valid = dataArb_io_out_valid;
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr;
  assign data_io_req_bits_write = dataArb_io_out_bits_write;
  assign data_io_req_bits_wdata = _T_124;
  assign data_io_req_bits_eccMask = dataArb_io_out_bits_eccMask;
  assign dataArb_io_in_0_valid = _T_1373;
  assign dataArb_io_in_0_bits_addr = _T_1453[13:0];
  assign dataArb_io_in_0_bits_write = 1'h1;
  assign dataArb_io_in_0_bits_wdata = _T_1455;
  assign dataArb_io_in_0_bits_eccMask = _T_1475;
  assign dataArb_io_in_1_valid = _GEN_122;
  assign dataArb_io_in_1_bits_addr = _T_3271[13:0];
  assign dataArb_io_in_1_bits_write = _GEN_123;
  assign dataArb_io_in_1_bits_wdata = io_mem_0_d_bits_data;
  assign dataArb_io_in_1_bits_eccMask = 4'hf;
  assign dataArb_io_in_2_valid = _T_3640;
  assign dataArb_io_in_2_bits_addr = _T_3644[13:0];
  assign dataArb_io_in_2_bits_write = 1'h0;
  assign dataArb_io_in_2_bits_wdata = 32'h0;
  assign dataArb_io_in_2_bits_eccMask = 4'h0;
  assign dataArb_io_in_3_valid = _T_356;
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[13:0];
  assign dataArb_io_in_3_bits_write = 1'h0;
  assign dataArb_io_in_3_bits_wdata = 32'h0;
  assign dataArb_io_in_3_bits_eccMask = 4'h0;
  assign dataArb_io_out_ready = 1'h1;
  assign _T_117 = dataArb_io_out_bits_wdata;
  assign _T_118 = _T_117[7:0];
  assign _T_119 = _T_117[15:8];
  assign _T_120 = _T_117[23:16];
  assign _T_121 = _T_117[31:24];
  assign _T_122 = {_T_119,_T_118};
  assign _T_123 = {_T_121,_T_120};
  assign _T_124 = {_T_123,_T_122};
  assign _T_133 = io_cpu_req_ready & io_cpu_req_valid;
  assign _T_136 = io_mem_0_b_ready & io_mem_0_b_valid;
  assign _GEN_2 = _T_136 ? io_mem_0_b_bits_param : probe_bits_param;
  assign _GEN_5 = _T_136 ? io_mem_0_b_bits_address : probe_bits_address;
  assign _T_144 = io_cpu_s1_kill == 1'h0;
  assign s1_valid_masked = s1_valid & _T_144;
  assign _T_146 = _GEN_152 == 1'h0;
  assign s1_valid_not_nacked = s1_valid & _T_146;
  assign _T_148 = metaArb_io_out_bits_write == 1'h0;
  assign _T_149 = metaArb_io_out_valid & _T_148;
  assign _T_150 = io_cpu_req_bits_addr[31:14];
  assign _T_151 = io_cpu_req_bits_addr[5:0];
  assign _T_152 = {_T_150,metaArb_io_out_bits_idx};
  assign _T_153 = {_T_152,_T_151};
  assign _GEN_8 = _T_149 ? _T_153 : s1_req_addr;
  assign _GEN_9 = _T_149 ? io_cpu_req_bits_tag : s1_req_tag;
  assign _GEN_10 = _T_149 ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign _GEN_11 = _T_149 ? io_cpu_req_bits_typ : s1_req_typ;
  assign _GEN_12 = _T_149 ? io_cpu_req_bits_phys : s1_req_phys;
  assign _T_155 = s1_req_cmd == 5'h0;
  assign _T_157 = s1_req_cmd == 5'h6;
  assign _T_158 = _T_155 | _T_157;
  assign _T_160 = s1_req_cmd == 5'h7;
  assign _T_161 = _T_158 | _T_160;
  assign _T_166 = s1_req_cmd == 5'h4;
  assign _T_167 = s1_req_cmd == 5'h9;
  assign _T_168 = s1_req_cmd == 5'ha;
  assign _T_169 = s1_req_cmd == 5'hb;
  assign _T_170 = _T_166 | _T_167;
  assign _T_171 = _T_170 | _T_168;
  assign _T_172 = _T_171 | _T_169;
  assign _T_178 = s1_req_cmd == 5'h8;
  assign _T_179 = s1_req_cmd == 5'hc;
  assign _T_180 = s1_req_cmd == 5'hd;
  assign _T_181 = s1_req_cmd == 5'he;
  assign _T_182 = s1_req_cmd == 5'hf;
  assign _T_183 = _T_178 | _T_179;
  assign _T_184 = _T_183 | _T_180;
  assign _T_185 = _T_184 | _T_181;
  assign _T_186 = _T_185 | _T_182;
  assign _T_187 = _T_172 | _T_186;
  assign s1_read = _T_161 | _T_187;
  assign _T_189 = s1_req_cmd == 5'h1;
  assign _T_191 = s1_req_cmd == 5'h11;
  assign _T_192 = _T_189 | _T_191;
  assign _T_195 = _T_192 | _T_160;
  assign s1_write = _T_195 | _T_187;
  assign s1_readwrite = s1_read | s1_write;
  assign s1_sfence = s1_req_cmd == 5'h14;
  assign _T_232 = release_state == 3'h1;
  assign _T_233 = release_state == 3'h2;
  assign inWriteback = _T_232 | _T_233;
  assign _T_235 = release_state == 3'h0;
  assign _T_237 = cached_grant_wait == 1'h0;
  assign _T_238 = _T_235 & _T_237;
  assign _T_241 = _T_238 & _T_146;
  assign _T_246 = io_cpu_req_bits_cmd == 5'h0;
  assign _T_248 = io_cpu_req_bits_cmd == 5'h6;
  assign _T_249 = _T_246 | _T_248;
  assign _T_251 = io_cpu_req_bits_cmd == 5'h7;
  assign _T_252 = _T_249 | _T_251;
  assign _T_257 = io_cpu_req_bits_cmd == 5'h4;
  assign _T_258 = io_cpu_req_bits_cmd == 5'h9;
  assign _T_259 = io_cpu_req_bits_cmd == 5'ha;
  assign _T_260 = io_cpu_req_bits_cmd == 5'hb;
  assign _T_261 = _T_257 | _T_258;
  assign _T_262 = _T_261 | _T_259;
  assign _T_263 = _T_262 | _T_260;
  assign _T_269 = io_cpu_req_bits_cmd == 5'h8;
  assign _T_270 = io_cpu_req_bits_cmd == 5'hc;
  assign _T_271 = io_cpu_req_bits_cmd == 5'hd;
  assign _T_272 = io_cpu_req_bits_cmd == 5'he;
  assign _T_273 = io_cpu_req_bits_cmd == 5'hf;
  assign _T_274 = _T_269 | _T_270;
  assign _T_275 = _T_274 | _T_271;
  assign _T_276 = _T_275 | _T_272;
  assign _T_277 = _T_276 | _T_273;
  assign _T_278 = _T_263 | _T_277;
  assign _T_279 = _T_252 | _T_278;
  assign _T_281 = io_cpu_req_bits_cmd == 5'h1;
  assign _T_283 = io_cpu_req_bits_cmd == 5'h11;
  assign _T_284 = _T_281 | _T_283;
  assign _T_287 = _T_284 | _T_251;
  assign _T_314 = _T_287 | _T_278;
  assign _T_321 = _T_314 & _T_283;
  assign s0_needsRead = _T_279 | _T_321;
  assign _T_356 = io_cpu_req_valid & s0_needsRead;
  assign _T_360 = 2'h1 << 1'h0;
  assign _T_364 = dataArb_io_in_3_ready == 1'h0;
  assign _T_365 = _T_364 & _T_279;
  assign _GEN_14 = _T_365 ? 1'h0 : _T_241;
  assign _T_375 = io_cpu_req_bits_addr[13:6];
  assign _T_379 = metaArb_io_in_7_ready == 1'h0;
  assign _GEN_16 = _T_379 ? 1'h0 : _GEN_14;
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = _T_385;
  assign tlb_io_req_bits_vaddr = s1_req_addr;
  assign tlb_io_req_bits_instruction = 1'h0;
  assign tlb_io_req_bits_size = s1_req_typ[1:0];
  assign tlb_io_req_bits_cmd = s1_req_cmd;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_sum = io_ptw_status_sum;
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr;
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask;
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr;
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask;
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr;
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask;
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr;
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask;
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr;
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask;
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr;
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask;
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr;
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask;
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr;
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask;
  assign _T_384 = s1_readwrite | s1_sfence;
  assign _T_385 = s1_valid_masked & _T_384;
  assign _T_390 = tlb_io_req_ready == 1'h0;
  assign _T_392 = tlb_io_ptw_resp_valid == 1'h0;
  assign _T_393 = _T_390 & _T_392;
  assign _T_395 = io_cpu_req_bits_phys == 1'h0;
  assign _T_396 = _T_393 & _T_395;
  assign _GEN_17 = _T_396 ? 1'h0 : _GEN_16;
  assign _T_398 = s1_valid & s1_readwrite;
  assign _T_399 = _T_398 & tlb_io_resp_miss;
  assign _T_408 = tlb_io_resp_paddr >= 32'h80000000;
  assign _T_410 = 32'h80000000 + 32'h4000;
  assign _T_411 = _T_410[31:0];
  assign _T_412 = tlb_io_resp_paddr < _T_411;
  assign s1_hit_way = _T_408 & _T_412;
  assign s1_hit_state_state = s1_hit_way ? 2'h3 : 2'h0;
  assign _T_428 = s1_req_typ[1:0];
  assign _T_430 = s1_req_addr[0];
  assign _T_434 = _T_428 >= 2'h1;
  assign _T_438 = _T_430 | _T_434;
  assign _T_441 = _T_430 ? 1'h0 : 1'h1;
  assign _T_442 = {_T_438,_T_441};
  assign _T_443 = s1_req_addr[1];
  assign _T_445 = _T_443 ? _T_442 : 2'h0;
  assign _T_447 = _T_428 >= 2'h2;
  assign _T_450 = _T_447 ? 2'h3 : 2'h0;
  assign _T_451 = _T_445 | _T_450;
  assign _T_454 = _T_443 ? 2'h0 : _T_442;
  assign _T_455 = {_T_451,_T_454};
  assign s1_mask = _T_191 ? io_cpu_s1_data_mask : _T_455;
  assign _T_457 = s1_sfence == 1'h0;
  assign _T_458 = s1_valid_masked & _T_457;
  assign _T_462 = {io_cpu_s2_xcpt_pf_st,io_cpu_s2_xcpt_ae_ld};
  assign _T_463 = {_T_462,io_cpu_s2_xcpt_ae_st};
  assign _T_464 = {io_cpu_s2_xcpt_ma_ld,io_cpu_s2_xcpt_ma_st};
  assign _T_465 = {_T_464,io_cpu_s2_xcpt_pf_ld};
  assign _T_466 = {_T_465,_T_463};
  assign _T_468 = _T_466 != 6'h0;
  assign _T_470 = _T_468 == 1'h0;
  assign s2_valid = _T_461 & _T_470;
  assign _T_473 = s1_probe | s2_probe;
  assign _T_474 = release_state != 3'h0;
  assign releaseInFlight = _T_473 | _T_474;
  assign s2_valid_masked = s2_valid & _T_478;
  assign _T_479 = s2_req_addr[31:6];
  assign _GEN_234 = {{6'd0}, _T_479};
  assign acquire_address = _GEN_234 << 6;
  assign _T_482 = s1_valid_not_nacked | s1_flush_valid;
  assign _GEN_19 = _T_482 ? tlb_io_resp_paddr : s2_req_addr;
  assign _GEN_20 = _T_482 ? s1_req_tag : s2_req_tag;
  assign _GEN_21 = _T_482 ? s1_req_cmd : s2_req_cmd;
  assign _GEN_22 = _T_482 ? s1_req_typ : s2_req_typ;
  assign _GEN_23 = _T_482 ? s1_req_phys : s2_req_phys;
  assign _GEN_25 = _T_482 ? 1'h1 : s2_uncached;
  assign _T_488 = s2_req_cmd == 5'h0;
  assign _T_490 = s2_req_cmd == 5'h6;
  assign _T_491 = _T_488 | _T_490;
  assign _T_493 = s2_req_cmd == 5'h7;
  assign _T_494 = _T_491 | _T_493;
  assign _T_499 = s2_req_cmd == 5'h4;
  assign _T_500 = s2_req_cmd == 5'h9;
  assign _T_501 = s2_req_cmd == 5'ha;
  assign _T_502 = s2_req_cmd == 5'hb;
  assign _T_503 = _T_499 | _T_500;
  assign _T_504 = _T_503 | _T_501;
  assign _T_505 = _T_504 | _T_502;
  assign _T_511 = s2_req_cmd == 5'h8;
  assign _T_512 = s2_req_cmd == 5'hc;
  assign _T_513 = s2_req_cmd == 5'hd;
  assign _T_514 = s2_req_cmd == 5'he;
  assign _T_515 = s2_req_cmd == 5'hf;
  assign _T_516 = _T_511 | _T_512;
  assign _T_517 = _T_516 | _T_513;
  assign _T_518 = _T_517 | _T_514;
  assign _T_519 = _T_518 | _T_515;
  assign _T_520 = _T_505 | _T_519;
  assign s2_read = _T_494 | _T_520;
  assign _T_522 = s2_req_cmd == 5'h1;
  assign _T_524 = s2_req_cmd == 5'h11;
  assign _T_525 = _T_522 | _T_524;
  assign _T_528 = _T_525 | _T_493;
  assign s2_write = _T_528 | _T_520;
  assign s2_readwrite = s2_read | s2_write;
  assign _T_571 = s1_valid | inWriteback;
  assign _GEN_27 = _T_571 ? data_io_resp_0 : s2_data;
  assign _GEN_29 = s1_probe ? s1_hit_state_state : s2_probe_state_state;
  assign _GEN_31 = s1_valid_not_nacked ? s1_hit_state_state : s2_hit_state_state;
  assign _GEN_32 = s1_valid_not_nacked ? 1'h0 : s2_waw_hazard;
  assign s2_hit_valid = s2_hit_state_state > 2'h0;
  assign _T_651 = s2_req_cmd == 5'h3;
  assign _T_652 = s2_write | _T_651;
  assign _T_655 = _T_652 | _T_490;
  assign _T_656 = {s2_write,_T_655};
  assign _T_657 = {_T_656,s2_hit_state_state};
  assign _T_744 = 4'hc == _T_657;
  assign _T_746 = _T_744 ? 2'h1 : 2'h0;
  assign _T_747 = 4'hd == _T_657;
  assign _T_749 = _T_747 ? 2'h2 : _T_746;
  assign _T_750 = 4'h4 == _T_657;
  assign _T_752 = _T_750 ? 2'h1 : _T_749;
  assign _T_753 = 4'h5 == _T_657;
  assign _T_755 = _T_753 ? 2'h2 : _T_752;
  assign _T_756 = 4'h0 == _T_657;
  assign _T_758 = _T_756 ? 2'h0 : _T_755;
  assign _T_759 = 4'he == _T_657;
  assign _T_761 = _T_759 ? 2'h3 : _T_758;
  assign _T_762 = 4'hf == _T_657;
  assign _T_763 = _T_762 ? 1'h1 : _T_759;
  assign _T_764 = _T_762 ? 2'h3 : _T_761;
  assign _T_765 = 4'h6 == _T_657;
  assign _T_766 = _T_765 ? 1'h1 : _T_763;
  assign _T_767 = _T_765 ? 2'h2 : _T_764;
  assign _T_768 = 4'h7 == _T_657;
  assign _T_769 = _T_768 ? 1'h1 : _T_766;
  assign _T_770 = _T_768 ? 2'h3 : _T_767;
  assign _T_771 = 4'h1 == _T_657;
  assign _T_772 = _T_771 ? 1'h1 : _T_769;
  assign _T_773 = _T_771 ? 2'h1 : _T_770;
  assign _T_774 = 4'h2 == _T_657;
  assign _T_775 = _T_774 ? 1'h1 : _T_772;
  assign _T_776 = _T_774 ? 2'h2 : _T_773;
  assign _T_777 = 4'h3 == _T_657;
  assign s2_hit = _T_777 ? 1'h1 : _T_775;
  assign s2_grow_param = _T_777 ? 2'h3 : _T_776;
  assign _T_779 = s2_data[7:0];
  assign _T_780 = s2_data[15:8];
  assign _T_781 = s2_data[23:16];
  assign _T_782 = s2_data[31:24];
  assign _T_855 = s2_req_typ[1:0];
  assign _T_876 = {_T_780,_T_779};
  assign _T_877 = {_T_782,_T_781};
  assign s2_data_corrected = {_T_877,_T_876};
  assign _T_880 = s2_valid_masked & s2_readwrite;
  assign s2_valid_hit_pre_data_ecc = _T_880 & s2_hit;
  assign _T_888 = s2_waw_hazard == 1'h0;
  assign s2_valid_hit = s2_valid_hit_pre_data_ecc & _T_888;
  assign _T_895 = s2_hit == 1'h0;
  assign _T_896 = _T_880 & _T_895;
  assign _T_898 = release_ack_wait == 1'h0;
  assign s2_valid_miss = _T_896 & _T_898;
  assign _T_900 = s2_uncached == 1'h0;
  assign _T_901 = s2_valid_miss & _T_900;
  assign _T_905 = uncachedInFlight_0 == 1'h0;
  assign s2_valid_cached_miss = _T_901 & _T_905;
  assign s2_valid_uncached = s2_valid_miss & s2_uncached;
  assign _T_910 = s2_flush_valid_pre_tag_ecc == 1'h0;
  assign _T_911 = s2_hit_valid & _T_910;
  assign _GEN_35 = _T_482 ? 2'h0 : _T_926_state;
  assign s2_victim_state_state = _T_911 ? s2_hit_state_state : _T_926_state;
  assign _T_927 = {probe_bits_param,s2_probe_state_state};
  assign _T_1015 = 4'hb == _T_927;
  assign _T_1019 = 4'h4 == _T_927;
  assign _T_1020 = _T_1019 ? 1'h0 : _T_1015;
  assign _T_1023 = 4'h5 == _T_927;
  assign _T_1024 = _T_1023 ? 1'h0 : _T_1020;
  assign _T_1027 = 4'h6 == _T_927;
  assign _T_1028 = _T_1027 ? 1'h0 : _T_1024;
  assign _T_1031 = 4'h7 == _T_927;
  assign _T_1032 = _T_1031 ? 1'h1 : _T_1028;
  assign _T_1035 = 4'h0 == _T_927;
  assign _T_1036 = _T_1035 ? 1'h0 : _T_1032;
  assign _T_1039 = 4'h1 == _T_927;
  assign _T_1040 = _T_1039 ? 1'h0 : _T_1036;
  assign _T_1043 = 4'h2 == _T_927;
  assign _T_1044 = _T_1043 ? 1'h0 : _T_1040;
  assign _T_1047 = 4'h3 == _T_927;
  assign s2_prb_ack_data = _T_1047 ? 1'h1 : _T_1044;
  assign _T_1064 = {2'h2,s2_victim_state_state};
  assign _T_1152 = 4'hb == _T_1064;
  assign _T_1156 = 4'h4 == _T_1064;
  assign _T_1157 = _T_1156 ? 1'h0 : _T_1152;
  assign _T_1160 = 4'h5 == _T_1064;
  assign _T_1161 = _T_1160 ? 1'h0 : _T_1157;
  assign _T_1164 = 4'h6 == _T_1064;
  assign _T_1165 = _T_1164 ? 1'h0 : _T_1161;
  assign _T_1168 = 4'h7 == _T_1064;
  assign _T_1169 = _T_1168 ? 1'h1 : _T_1165;
  assign _T_1172 = 4'h0 == _T_1064;
  assign _T_1173 = _T_1172 ? 1'h0 : _T_1169;
  assign _T_1176 = 4'h1 == _T_1064;
  assign _T_1177 = _T_1176 ? 1'h0 : _T_1173;
  assign _T_1180 = 4'h2 == _T_1064;
  assign _T_1181 = _T_1180 ? 1'h0 : _T_1177;
  assign _T_1184 = 4'h3 == _T_1064;
  assign s2_victim_dirty = _T_1184 ? 1'h1 : _T_1181;
  assign _T_1187 = s2_hit_state_state == s2_grow_param;
  assign s2_update_meta = _T_1187 == 1'h0;
  assign _T_1190 = s2_valid_hit == 1'h0;
  assign _T_1191 = s2_valid & _T_1190;
  assign _T_1192 = s2_valid_uncached & io_mem_0_a_ready;
  assign _T_1193 = ~ uncachedInFlight_0;
  assign _T_1195 = _T_1193 == 1'h0;
  assign _T_1197 = _T_1195 == 1'h0;
  assign _T_1198 = _T_1192 & _T_1197;
  assign _T_1200 = _T_1198 == 1'h0;
  assign _T_1201 = _T_1191 & _T_1200;
  assign _T_1202 = s2_valid_hit & s2_update_meta;
  assign _T_1203 = io_cpu_s2_nack | _T_1202;
  assign _GEN_36 = _T_1203 ? 1'h1 : _T_399;
  assign _T_1214 = s2_probe ? probe_bits_address : s2_req_addr;
  assign _T_1215 = _T_1214[13:6];
  assign _T_1219 = s2_victim_dirty == 1'h0;
  assign _T_1223 = s2_req_addr[13:6];
  assign lrscValid = lrscCount > 5'h3;
  assign _T_1248 = lrscCount > 5'h0;
  assign _T_1250 = lrscCount - 5'h1;
  assign _T_1251 = $unsigned(_T_1250);
  assign _T_1252 = _T_1251[4:0];
  assign _GEN_39 = _T_1248 ? _T_1252 : lrscCount;
  assign _T_1255 = s2_valid_masked & _T_1248;
  assign _T_1256 = _T_1255 | io_cpu_invalidate_lr;
  assign _GEN_40 = _T_1256 ? 5'h0 : _GEN_39;
  assign _T_1262 = s1_valid_not_nacked & s1_write;
  assign _GEN_41 = _T_1262 ? s1_req_cmd : pstore1_cmd;
  assign _GEN_42 = _T_1262 ? tlb_io_resp_paddr : pstore1_addr;
  assign _GEN_43 = _T_1262 ? io_cpu_s1_data_data : a_data;
  assign _GEN_45 = _T_1262 ? s1_mask : pstore1_mask;
  assign _T_1350 = s1_write & _T_191;
  assign _T_1351 = s1_read | _T_1350;
  assign _GEN_46 = _T_1262 ? _T_1351 : _T_1354;
  assign _T_1358 = _T_1396 & pstore2_valid;
  assign _T_1359 = s1_valid & s1_write;
  assign _T_1360 = _T_1359 | _T_1354;
  assign pstore_drain_structural = _T_1358 & _T_1360;
  assign pstore_drain_opportunistic = _T_356 == 1'h0;
  assign pstore_drain_on_miss = releaseInFlight | io_cpu_s2_nack;
  assign _T_1368 = _T_1354 == 1'h0;
  assign _T_1369 = _T_1396 & _T_1368;
  assign _T_1370 = _T_1369 | pstore2_valid;
  assign _T_1371 = pstore_drain_opportunistic | pstore_drain_on_miss;
  assign _T_1372 = _T_1370 & _T_1371;
  assign _T_1373 = pstore_drain_structural | _T_1372;
  assign _T_1374 = s2_valid_hit & s2_write;
  assign _T_1381 = _T_1374 == 1'h0;
  assign _T_1383 = _T_1379 == 1'h0;
  assign _T_1384 = _T_1381 | _T_1383;
  assign _T_1385 = _T_1384 | reset;
  assign _T_1387 = _T_1385 == 1'h0;
  assign _T_1391 = _T_1374 | _T_1379;
  assign _T_1392 = _T_1391 & pstore2_valid;
  assign _T_1394 = _T_1373 == 1'h0;
  assign _T_1395 = _T_1392 & _T_1394;
  assign _T_1396 = _T_1374 | _T_1379;
  assign _T_1398 = pstore2_valid == _T_1373;
  assign advance_pstore1 = _T_1391 & _T_1398;
  assign _T_1401 = pstore2_valid & _T_1394;
  assign _T_1402 = _T_1401 | advance_pstore1;
  assign _GEN_47 = advance_pstore1 ? pstore1_addr : pstore2_addr;
  assign _T_1408 = pstore2_addr[13:2];
  assign _T_1417 = _GEN_216[7:0];
  assign _T_1418 = pstore1_mask[0];
  assign _GEN_49 = advance_pstore1 ? _T_1417 : _T_1422;
  assign _T_1423 = _GEN_216[15:8];
  assign _T_1424 = pstore1_mask[1];
  assign _GEN_50 = advance_pstore1 ? _T_1423 : _T_1428;
  assign _T_1429 = _GEN_216[23:16];
  assign _T_1430 = pstore1_mask[2];
  assign _GEN_51 = advance_pstore1 ? _T_1429 : _T_1434;
  assign _T_1435 = _GEN_216[31:24];
  assign _T_1436 = pstore1_mask[3];
  assign _GEN_52 = advance_pstore1 ? _T_1435 : _T_1440;
  assign _T_1441 = {_T_1428,_T_1422};
  assign _T_1442 = {_T_1440,_T_1434};
  assign pstore2_storegen_data = {_T_1442,_T_1441};
  assign _T_1449 = ~ pstore1_mask;
  assign _T_1451 = ~ _T_1449;
  assign _GEN_53 = advance_pstore1 ? _T_1451 : pstore2_storegen_mask;
  assign _T_1453 = pstore2_valid ? pstore2_addr : pstore1_addr;
  assign _T_1455 = pstore2_valid ? pstore2_storegen_data : a_data;
  assign _T_1460 = pstore2_valid ? pstore2_storegen_mask : pstore1_mask;
  assign _T_1461 = _T_1460[0];
  assign _T_1462 = _T_1460[1];
  assign _T_1463 = _T_1460[2];
  assign _T_1464 = _T_1460[3];
  assign _T_1473 = {_T_1462,_T_1461};
  assign _T_1474 = {_T_1464,_T_1463};
  assign _T_1475 = {_T_1474,_T_1473};
  assign _T_1476 = pstore1_addr[13:2];
  assign _T_1477 = s1_req_addr[13:2];
  assign _T_1478 = _T_1476 == _T_1477;
  assign _T_1491 = {_T_1424,_T_1418};
  assign _T_1492 = {_T_1436,_T_1430};
  assign _T_1493 = {_T_1492,_T_1491};
  assign _T_1494 = _T_1493[0];
  assign _T_1495 = _T_1493[1];
  assign _T_1496 = _T_1493[2];
  assign _T_1497 = _T_1493[3];
  assign _T_1498 = {_T_1495,_T_1494};
  assign _T_1499 = {_T_1497,_T_1496};
  assign _T_1500 = {_T_1499,_T_1498};
  assign _T_1501 = s1_mask[0];
  assign _T_1502 = s1_mask[1];
  assign _T_1503 = s1_mask[2];
  assign _T_1504 = s1_mask[3];
  assign _T_1513 = {_T_1502,_T_1501};
  assign _T_1514 = {_T_1504,_T_1503};
  assign _T_1515 = {_T_1514,_T_1513};
  assign _T_1516 = _T_1515[0];
  assign _T_1517 = _T_1515[1];
  assign _T_1518 = _T_1515[2];
  assign _T_1519 = _T_1515[3];
  assign _T_1520 = {_T_1517,_T_1516};
  assign _T_1521 = {_T_1519,_T_1518};
  assign _T_1522 = {_T_1521,_T_1520};
  assign _T_1523 = _T_1500 & _T_1522;
  assign _T_1525 = _T_1523 != 4'h0;
  assign _T_1526 = pstore1_mask & s1_mask;
  assign _T_1528 = _T_1526 != 4'h0;
  assign _T_1529 = s1_write ? _T_1525 : _T_1528;
  assign _T_1530 = _T_1478 & _T_1529;
  assign _T_1531 = _T_1391 & _T_1530;
  assign _T_1534 = _T_1408 == _T_1477;
  assign _T_1535 = pstore2_storegen_mask[0];
  assign _T_1536 = pstore2_storegen_mask[1];
  assign _T_1537 = pstore2_storegen_mask[2];
  assign _T_1538 = pstore2_storegen_mask[3];
  assign _T_1547 = {_T_1536,_T_1535};
  assign _T_1548 = {_T_1538,_T_1537};
  assign _T_1549 = {_T_1548,_T_1547};
  assign _T_1550 = _T_1549[0];
  assign _T_1551 = _T_1549[1];
  assign _T_1552 = _T_1549[2];
  assign _T_1553 = _T_1549[3];
  assign _T_1554 = {_T_1551,_T_1550};
  assign _T_1555 = {_T_1553,_T_1552};
  assign _T_1556 = {_T_1555,_T_1554};
  assign _T_1579 = _T_1556 & _T_1522;
  assign _T_1581 = _T_1579 != 4'h0;
  assign _T_1582 = pstore2_storegen_mask & s1_mask;
  assign _T_1584 = _T_1582 != 4'h0;
  assign _T_1585 = s1_write ? _T_1581 : _T_1584;
  assign _T_1586 = _T_1534 & _T_1585;
  assign _T_1587 = pstore2_valid & _T_1586;
  assign s1_hazard = _T_1531 | _T_1587;
  assign s1_raw_hazard = s1_read & s1_hazard;
  assign _T_1592 = s1_valid & s1_raw_hazard;
  assign _GEN_54 = _T_1592 ? 1'h1 : _GEN_36;
  assign acquire__param = {{1'd0}, s2_grow_param};
  assign get_size = {{2'd0}, _T_855};
  assign _T_1799 = _T_855[0];
  assign _T_1801 = 2'h1 << _T_1799;
  assign _T_1804 = _T_1801 | 2'h1;
  assign _T_1806 = _T_855 >= 2'h2;
  assign _T_1808 = _T_1804[1];
  assign _T_1809 = s2_req_addr[1];
  assign _T_1811 = _T_1809 == 1'h0;
  assign _T_1813 = _T_1808 & _T_1811;
  assign _T_1814 = _T_1806 | _T_1813;
  assign _T_1816 = _T_1808 & _T_1809;
  assign _T_1817 = _T_1806 | _T_1816;
  assign _T_1818 = _T_1804[0];
  assign _T_1819 = s2_req_addr[0];
  assign _T_1821 = _T_1819 == 1'h0;
  assign _T_1822 = _T_1811 & _T_1821;
  assign _T_1823 = _T_1818 & _T_1822;
  assign _T_1824 = _T_1814 | _T_1823;
  assign _T_1825 = _T_1811 & _T_1819;
  assign _T_1826 = _T_1818 & _T_1825;
  assign _T_1827 = _T_1814 | _T_1826;
  assign _T_1828 = _T_1809 & _T_1821;
  assign _T_1829 = _T_1818 & _T_1828;
  assign _T_1830 = _T_1817 | _T_1829;
  assign _T_1831 = _T_1809 & _T_1819;
  assign _T_1832 = _T_1818 & _T_1831;
  assign _T_1833 = _T_1817 | _T_1832;
  assign _T_1834 = {_T_1827,_T_1824};
  assign _T_1835 = {_T_1833,_T_1830};
  assign _T_1836 = {_T_1835,_T_1834};
  assign put_size = {{2'd0}, _T_855};
  assign _T_2060_size = {{2'd0}, _T_855};
  assign _T_2187_size = {{2'd0}, _T_855};
  assign _T_2314_size = {{2'd0}, _T_855};
  assign _T_2441_size = {{2'd0}, _T_855};
  assign _T_2568_size = {{2'd0}, _T_855};
  assign _T_2695_size = {{2'd0}, _T_855};
  assign _T_2822_size = {{2'd0}, _T_855};
  assign _T_2949_size = {{2'd0}, _T_855};
  assign _T_3076_size = {{2'd0}, _T_855};
  assign _T_3116 = 5'hf == s2_req_cmd;
  assign _T_3117_opcode = _T_3116 ? 3'h2 : 3'h0;
  assign _T_3117_param = _T_3116 ? 3'h3 : 3'h0;
  assign _T_3117_size = _T_3116 ? _T_3076_size : 4'h0;
  assign _T_3117_address = _T_3116 ? s2_req_addr : 32'h0;
  assign _T_3117_mask = _T_3116 ? _T_1836 : 4'h0;
  assign _T_3117_data = _T_3116 ? a_data : 32'h0;
  assign _T_3118 = 5'he == s2_req_cmd;
  assign _T_3119_opcode = _T_3118 ? 3'h2 : _T_3117_opcode;
  assign _T_3119_param = _T_3118 ? 3'h2 : _T_3117_param;
  assign _T_3119_size = _T_3118 ? _T_2949_size : _T_3117_size;
  assign _T_3119_address = _T_3118 ? s2_req_addr : _T_3117_address;
  assign _T_3119_mask = _T_3118 ? _T_1836 : _T_3117_mask;
  assign _T_3119_data = _T_3118 ? a_data : _T_3117_data;
  assign _T_3120 = 5'hd == s2_req_cmd;
  assign _T_3121_opcode = _T_3120 ? 3'h2 : _T_3119_opcode;
  assign _T_3121_param = _T_3120 ? 3'h1 : _T_3119_param;
  assign _T_3121_size = _T_3120 ? _T_2822_size : _T_3119_size;
  assign _T_3121_address = _T_3120 ? s2_req_addr : _T_3119_address;
  assign _T_3121_mask = _T_3120 ? _T_1836 : _T_3119_mask;
  assign _T_3121_data = _T_3120 ? a_data : _T_3119_data;
  assign _T_3122 = 5'hc == s2_req_cmd;
  assign _T_3123_opcode = _T_3122 ? 3'h2 : _T_3121_opcode;
  assign _T_3123_param = _T_3122 ? 3'h0 : _T_3121_param;
  assign _T_3123_size = _T_3122 ? _T_2695_size : _T_3121_size;
  assign _T_3123_address = _T_3122 ? s2_req_addr : _T_3121_address;
  assign _T_3123_mask = _T_3122 ? _T_1836 : _T_3121_mask;
  assign _T_3123_data = _T_3122 ? a_data : _T_3121_data;
  assign _T_3124 = 5'h8 == s2_req_cmd;
  assign _T_3125_opcode = _T_3124 ? 3'h2 : _T_3123_opcode;
  assign _T_3125_param = _T_3124 ? 3'h4 : _T_3123_param;
  assign _T_3125_size = _T_3124 ? _T_2568_size : _T_3123_size;
  assign _T_3125_address = _T_3124 ? s2_req_addr : _T_3123_address;
  assign _T_3125_mask = _T_3124 ? _T_1836 : _T_3123_mask;
  assign _T_3125_data = _T_3124 ? a_data : _T_3123_data;
  assign _T_3126 = 5'hb == s2_req_cmd;
  assign _T_3127_opcode = _T_3126 ? 3'h3 : _T_3125_opcode;
  assign _T_3127_param = _T_3126 ? 3'h2 : _T_3125_param;
  assign _T_3127_size = _T_3126 ? _T_2441_size : _T_3125_size;
  assign _T_3127_address = _T_3126 ? s2_req_addr : _T_3125_address;
  assign _T_3127_mask = _T_3126 ? _T_1836 : _T_3125_mask;
  assign _T_3127_data = _T_3126 ? a_data : _T_3125_data;
  assign _T_3128 = 5'ha == s2_req_cmd;
  assign _T_3129_opcode = _T_3128 ? 3'h3 : _T_3127_opcode;
  assign _T_3129_param = _T_3128 ? 3'h1 : _T_3127_param;
  assign _T_3129_size = _T_3128 ? _T_2314_size : _T_3127_size;
  assign _T_3129_address = _T_3128 ? s2_req_addr : _T_3127_address;
  assign _T_3129_mask = _T_3128 ? _T_1836 : _T_3127_mask;
  assign _T_3129_data = _T_3128 ? a_data : _T_3127_data;
  assign _T_3130 = 5'h9 == s2_req_cmd;
  assign _T_3131_opcode = _T_3130 ? 3'h3 : _T_3129_opcode;
  assign _T_3131_param = _T_3130 ? 3'h0 : _T_3129_param;
  assign _T_3131_size = _T_3130 ? _T_2187_size : _T_3129_size;
  assign _T_3131_address = _T_3130 ? s2_req_addr : _T_3129_address;
  assign _T_3131_mask = _T_3130 ? _T_1836 : _T_3129_mask;
  assign _T_3131_data = _T_3130 ? a_data : _T_3129_data;
  assign _T_3132 = 5'h4 == s2_req_cmd;
  assign atomics_opcode = _T_3132 ? 3'h3 : _T_3131_opcode;
  assign atomics_param = _T_3132 ? 3'h3 : _T_3131_param;
  assign atomics_size = _T_3132 ? _T_2060_size : _T_3131_size;
  assign atomics_address = _T_3132 ? s2_req_addr : _T_3131_address;
  assign atomics_mask = _T_3132 ? _T_1836 : _T_3131_mask;
  assign atomics_data = _T_3132 ? a_data : _T_3131_data;
  assign _T_3137 = s2_valid_cached_miss & _T_1219;
  assign _T_3143 = s2_valid_uncached & _T_1197;
  assign _T_3144 = _T_3137 | _T_3143;
  assign _T_3148 = s2_write == 1'h0;
  assign _T_3150 = s2_read == 1'h0;
  assign _T_3151_opcode = _T_3150 ? 3'h0 : atomics_opcode;
  assign _T_3151_param = _T_3150 ? 3'h0 : atomics_param;
  assign _T_3151_size = _T_3150 ? put_size : atomics_size;
  assign _T_3151_address = _T_3150 ? s2_req_addr : atomics_address;
  assign _T_3151_mask = _T_3150 ? _T_1836 : atomics_mask;
  assign _T_3151_data = _T_3150 ? a_data : atomics_data;
  assign _T_3152_opcode = _T_3148 ? 3'h4 : _T_3151_opcode;
  assign _T_3152_param = _T_3148 ? 3'h0 : _T_3151_param;
  assign _T_3152_size = _T_3148 ? get_size : _T_3151_size;
  assign _T_3152_address = _T_3148 ? s2_req_addr : _T_3151_address;
  assign _T_3152_mask = _T_3148 ? _T_1836 : _T_3151_mask;
  assign _T_3152_data = _T_3148 ? 32'h0 : _T_3151_data;
  assign _T_3153_opcode = _T_900 ? 3'h6 : _T_3152_opcode;
  assign _T_3153_param = _T_900 ? acquire__param : _T_3152_param;
  assign _T_3153_size = _T_900 ? 4'h6 : _T_3152_size;
  assign _T_3153_address = _T_900 ? acquire_address : _T_3152_address;
  assign _T_3153_mask = _T_900 ? 4'hf : _T_3152_mask;
  assign _T_3153_data = _T_900 ? 32'h0 : _T_3152_data;
  assign _T_3157 = _T_360[0];
  assign _T_3158 = io_mem_0_a_ready & _T_3144;
  assign _GEN_55 = _T_3157 ? 1'h1 : uncachedInFlight_0;
  assign _GEN_56 = _T_3157 ? s2_req_addr : uncachedReqs_0_addr;
  assign _GEN_57 = _T_3157 ? s2_req_tag : uncachedReqs_0_tag;
  assign _GEN_59 = _T_3157 ? s2_req_typ : uncachedReqs_0_typ;
  assign _GEN_62 = s2_uncached ? _GEN_55 : uncachedInFlight_0;
  assign _GEN_63 = s2_uncached ? _GEN_56 : uncachedReqs_0_addr;
  assign _GEN_64 = s2_uncached ? _GEN_57 : uncachedReqs_0_tag;
  assign _GEN_66 = s2_uncached ? _GEN_59 : uncachedReqs_0_typ;
  assign _GEN_69 = _T_900 ? 1'h1 : cached_grant_wait;
  assign _GEN_70 = _T_3158 ? _GEN_62 : uncachedInFlight_0;
  assign _GEN_71 = _T_3158 ? _GEN_63 : uncachedReqs_0_addr;
  assign _GEN_72 = _T_3158 ? _GEN_64 : uncachedReqs_0_tag;
  assign _GEN_74 = _T_3158 ? _GEN_66 : uncachedReqs_0_typ;
  assign _GEN_77 = _T_3158 ? _GEN_69 : cached_grant_wait;
  assign _T_3164 = io_mem_0_d_ready & io_mem_0_d_valid;
  assign _T_3167 = 27'hfff << io_mem_0_d_bits_size;
  assign _T_3168 = _T_3167[11:0];
  assign _T_3169 = ~ _T_3168;
  assign _T_3170 = _T_3169[11:2];
  assign _T_3171 = io_mem_0_d_bits_opcode[0];
  assign _T_3173 = _T_3171 ? _T_3170 : 10'h0;
  assign _T_3178 = _T_3176 - 10'h1;
  assign _T_3179 = $unsigned(_T_3178);
  assign _T_3180 = _T_3179[9:0];
  assign d_first = _T_3176 == 10'h0;
  assign _T_3183 = _T_3176 == 10'h1;
  assign _T_3185 = _T_3173 == 10'h0;
  assign d_last = _T_3183 | _T_3185;
  assign d_done = d_last & _T_3164;
  assign _T_3186 = ~ _T_3180;
  assign _T_3187 = _T_3173 & _T_3186;
  assign _T_3188 = d_first ? _T_3173 : _T_3180;
  assign _GEN_78 = _T_3164 ? _T_3188 : _T_3176;
  assign _GEN_235 = {{2'd0}, _T_3187};
  assign d_address_inc = _GEN_235 << 2;
  assign _T_3191 = io_mem_0_d_bits_opcode == 3'h4;
  assign _T_3192 = io_mem_0_d_bits_opcode == 3'h5;
  assign grantIsCached = _T_3191 | _T_3192;
  assign _T_3196 = io_mem_0_d_bits_opcode == 3'h0;
  assign _T_3197 = io_mem_0_d_bits_opcode == 3'h1;
  assign _T_3198 = io_mem_0_d_bits_opcode == 3'h2;
  assign _T_3199 = _T_3196 | _T_3197;
  assign grantIsUncached = _T_3199 | _T_3198;
  assign grantIsVoluntary = io_mem_0_d_bits_opcode == 3'h6;
  assign _T_3208 = blockProbeAfterGrantCount > 3'h0;
  assign _T_3210 = blockProbeAfterGrantCount - 3'h1;
  assign _T_3211 = $unsigned(_T_3210);
  assign _T_3212 = _T_3211[2:0];
  assign _GEN_79 = _T_3208 ? _T_3212 : blockProbeAfterGrantCount;
  assign _T_3214 = d_first == 1'h0;
  assign _T_3215 = _T_3214 | io_mem_0_e_ready;
  assign _T_3218 = grantIsCached ? _T_3215 : 1'h1;
  assign _T_3221 = cached_grant_wait | reset;
  assign _T_3223 = _T_3221 == 1'h0;
  assign _GEN_80 = d_last ? 1'h0 : _GEN_77;
  assign _GEN_81 = d_last ? 1'h0 : 1'h1;
  assign _GEN_82 = d_last ? 3'h7 : _GEN_79;
  assign _GEN_84 = grantIsCached ? _GEN_81 : grantInProgress;
  assign _GEN_85 = grantIsCached ? _GEN_80 : _GEN_77;
  assign _GEN_86 = grantIsCached ? _GEN_82 : _GEN_79;
  assign _T_3229 = grantIsCached == 1'h0;
  assign _T_3230 = _T_3229 & grantIsUncached;
  assign _T_3233 = 2'h1 << io_mem_0_d_bits_source;
  assign _T_3234 = _T_3233[0];
  assign _T_3238 = _T_3234 & d_last;
  assign _T_3239 = uncachedInFlight_0 | reset;
  assign _T_3241 = _T_3239 == 1'h0;
  assign _GEN_88 = _T_3238 ? 1'h0 : _GEN_70;
  assign _T_3243 = io_mem_0_d_bits_data[7:0];
  assign _T_3244 = io_mem_0_d_bits_data[15:8];
  assign _T_3245 = io_mem_0_d_bits_data[23:16];
  assign _T_3246 = io_mem_0_d_bits_data[31:24];
  assign _T_3247 = {_T_3244,_T_3243};
  assign _T_3248 = {_T_3246,_T_3245};
  assign _T_3249 = {_T_3248,_T_3247};
  assign _T_3251 = tlb_io_resp_paddr[31:2];
  assign _T_3252 = uncachedReqs_0_addr[1:0];
  assign _T_3253 = {_T_3251,_T_3252};
  assign _GEN_89 = _T_3197 ? _T_3249 : _GEN_27;
  assign _GEN_90 = _T_3197 ? 5'h0 : _GEN_21;
  assign _GEN_91 = _T_3197 ? uncachedReqs_0_typ : _GEN_22;
  assign _GEN_92 = _T_3197 ? uncachedReqs_0_tag : _GEN_20;
  assign _GEN_93 = _T_3197 ? _T_3253 : _GEN_19;
  assign _GEN_95 = _T_3230 ? _GEN_88 : _GEN_70;
  assign _GEN_96 = _T_3230 ? _GEN_89 : _GEN_27;
  assign _GEN_97 = _T_3230 ? _GEN_90 : _GEN_21;
  assign _GEN_98 = _T_3230 ? _GEN_91 : _GEN_22;
  assign _GEN_99 = _T_3230 ? _GEN_92 : _GEN_20;
  assign _GEN_100 = _T_3230 ? _GEN_93 : _GEN_19;
  assign _T_3257 = grantIsUncached == 1'h0;
  assign _T_3258 = _T_3229 & _T_3257;
  assign _T_3259 = _T_3258 & grantIsVoluntary;
  assign _T_3260 = release_ack_wait | reset;
  assign _T_3262 = _T_3260 == 1'h0;
  assign _GEN_102 = _T_3259 ? 1'h0 : release_ack_wait;
  assign _GEN_103 = _T_3164 ? _GEN_84 : grantInProgress;
  assign _GEN_104 = _T_3164 ? _GEN_85 : _GEN_77;
  assign _GEN_105 = _T_3164 ? _GEN_86 : _GEN_79;
  assign _GEN_107 = _T_3164 ? _GEN_95 : _GEN_70;
  assign _GEN_108 = _T_3164 ? _GEN_96 : _GEN_27;
  assign _GEN_109 = _T_3164 ? _GEN_97 : _GEN_21;
  assign _GEN_110 = _T_3164 ? _GEN_98 : _GEN_22;
  assign _GEN_111 = _T_3164 ? _GEN_99 : _GEN_20;
  assign _GEN_112 = _T_3164 ? _GEN_100 : _GEN_19;
  assign _GEN_114 = _T_3164 ? _GEN_102 : release_ack_wait;
  assign _T_3264 = io_mem_0_d_valid & _T_3192;
  assign _T_3267 = dataArb_io_in_1_ready == 1'h0;
  assign _T_3268 = _T_3192 & _T_3267;
  assign _GEN_115 = _T_3268 ? 1'h0 : _T_3218;
  assign _GEN_236 = {{20'd0}, d_address_inc};
  assign _T_3271 = acquire_address | _GEN_236;
  assign _T_3276 = grantIsCached & d_done;
  assign _T_3278 = metaArb_io_in_3_valid == 1'h0;
  assign _T_3279 = _T_3278 | metaArb_io_in_3_ready;
  assign _T_3280 = _T_3279 | reset;
  assign _T_3282 = _T_3280 == 1'h0;
  assign _T_3400 = blockUncachedGrant | s1_valid;
  assign _T_3401 = _T_3197 & _T_3400;
  assign _GEN_116 = io_mem_0_d_valid ? 1'h0 : _GEN_17;
  assign _GEN_117 = io_mem_0_d_valid ? 1'h1 : _T_3264;
  assign _GEN_118 = io_mem_0_d_valid ? 1'h0 : 1'h1;
  assign _GEN_119 = io_mem_0_d_valid ? _T_3267 : dataArb_io_out_valid;
  assign _GEN_120 = _T_3401 ? 1'h0 : _GEN_115;
  assign _GEN_121 = _T_3401 ? _GEN_116 : _GEN_17;
  assign _GEN_122 = _T_3401 ? _GEN_117 : _T_3264;
  assign _GEN_123 = _T_3401 ? _GEN_118 : 1'h1;
  assign _GEN_124 = _T_3401 ? _GEN_119 : dataArb_io_out_valid;
  assign _T_3408 = io_mem_0_d_valid & d_first;
  assign _T_3409 = _T_3408 & grantIsCached;
  assign _T_3413 = io_mem_0_e_ready & io_mem_0_e_valid;
  assign _T_3415 = _T_3164 | reset;
  assign _T_3417 = _T_3415 == 1'h0;
  assign _T_3418 = releaseInFlight | grantInProgress;
  assign _T_3421 = _T_3418 | _T_3208;
  assign _T_3422 = _T_3421 | lrscValid;
  assign _T_3425 = _T_3422 == 1'h0;
  assign _T_3426 = io_mem_0_b_valid & _T_3425;
  assign _T_3429 = metaArb_io_in_6_ready & _T_3425;
  assign _T_3431 = s1_valid == 1'h0;
  assign _T_3432 = _T_3429 & _T_3431;
  assign _T_3434 = s2_valid == 1'h0;
  assign _T_3435 = _T_3434 | s2_valid_hit;
  assign _T_3436 = _T_3432 & _T_3435;
  assign _T_3438 = io_mem_0_b_bits_address[13:6];
  assign _T_3441 = io_mem_0_c_ready & io_mem_0_c_valid;
  assign _T_3456 = _T_3454 - 10'h1;
  assign _T_3457 = $unsigned(_T_3456);
  assign _T_3458 = _T_3457[9:0];
  assign c_first = _T_3454 == 10'h0;
  assign _T_3465 = c_first ? 10'h0 : _T_3458;
  assign _GEN_125 = _T_3441 ? _T_3465 : _T_3454;
  assign _T_3467 = io_mem_0_c_ready == 1'h0;
  assign releaseRejected = io_mem_0_c_valid & _T_3467;
  assign _T_3468 = dataArb_io_in_2_ready & dataArb_io_in_2_valid;
  assign _T_3471 = releaseRejected == 1'h0;
  assign _T_3472 = s1_release_data_valid & _T_3471;
  assign _T_3478 = {1'h0,s2_release_data_valid};
  assign _GEN_237 = {{1'd0}, s1_release_data_valid};
  assign _T_3479 = _GEN_237 + _T_3478;
  assign _T_3480 = _T_3479[1:0];
  assign _T_3481 = releaseRejected ? 2'h0 : _T_3480;
  assign _GEN_238 = {{9'd0}, _T_3481};
  assign _T_3482 = 11'h0 + _GEN_238;
  assign releaseDataBeat = _T_3482[10:0];
  assign _GEN_129 = s2_prb_ack_data ? 3'h2 : release_state;
  assign _T_3517 = s2_probe_state_state > 2'h0;
  assign _T_3521 = s2_prb_ack_data == 1'h0;
  assign _T_3523 = _T_3521 & _T_3517;
  assign _T_3525 = _T_3441 ? 3'h7 : 3'h3;
  assign _GEN_130 = _T_3523 ? 1'h1 : s2_release_data_valid;
  assign _GEN_138 = _T_3523 ? _T_3525 : _GEN_129;
  assign _T_3532 = _T_3517 == 1'h0;
  assign _T_3533 = _T_3521 & _T_3532;
  assign _T_3536 = _T_3441 == 1'h0;
  assign _T_3537 = _T_3441 ? 3'h0 : 3'h5;
  assign _GEN_139 = _T_3533 ? 1'h1 : _GEN_130;
  assign _GEN_140 = _T_3533 ? _T_3536 : 1'h1;
  assign _GEN_141 = _T_3533 ? _T_3537 : _GEN_138;
  assign _GEN_142 = _GEN_140 ? 1'h1 : _GEN_54;
  assign _GEN_143 = s2_probe ? _GEN_141 : release_state;
  assign _GEN_144 = s2_probe ? _GEN_139 : s2_release_data_valid;
  assign _GEN_152 = s2_probe ? _GEN_142 : _GEN_54;
  assign _T_3539 = release_state == 3'h4;
  assign _T_3541 = probe_bits_address[13:6];
  assign _GEN_153 = metaArb_io_in_6_ready ? 3'h0 : _GEN_143;
  assign _GEN_154 = metaArb_io_in_6_ready ? 1'h1 : _T_136;
  assign _GEN_155 = _T_3539 ? 1'h1 : _T_3426;
  assign _GEN_156 = _T_3539 ? _T_3541 : _T_3438;
  assign _GEN_157 = _T_3539 ? _GEN_153 : _GEN_143;
  assign _GEN_158 = _T_3539 ? _GEN_154 : _T_136;
  assign _T_3543 = release_state == 3'h5;
  assign _GEN_159 = _T_3441 ? 3'h0 : _GEN_157;
  assign _GEN_160 = _T_3543 ? 1'h1 : _GEN_144;
  assign _GEN_161 = _T_3543 ? _GEN_159 : _GEN_157;
  assign _T_3545 = release_state == 3'h3;
  assign _GEN_162 = _T_3441 ? 3'h7 : _GEN_161;
  assign _GEN_163 = _T_3545 ? 1'h1 : _GEN_160;
  assign _GEN_171 = _T_3545 ? _GEN_162 : _GEN_161;
  assign _GEN_172 = _T_3441 ? 3'h7 : _GEN_171;
  assign _GEN_180 = _T_233 ? _GEN_172 : _GEN_171;
  assign _T_3549 = release_state == 3'h6;
  assign _T_3550 = _T_232 | _T_3549;
  assign _GEN_181 = _T_3441 ? 3'h6 : _GEN_180;
  assign _T_3636 = _T_3441 & c_first;
  assign _GEN_182 = _T_3636 ? 1'h1 : _GEN_114;
  assign _GEN_192 = _T_3550 ? _GEN_181 : _GEN_180;
  assign _GEN_193 = _T_3550 ? _GEN_182 : _GEN_114;
  assign _T_3639 = releaseDataBeat < 11'h10;
  assign _T_3640 = inWriteback & _T_3639;
  assign _T_3642 = releaseDataBeat[3:0];
  assign _GEN_246 = {{2'd0}, _T_3642};
  assign _T_3643 = _GEN_246 << 2;
  assign _GEN_247 = {{26'd0}, _T_3643};
  assign _T_3644 = io_mem_0_c_bits_address | _GEN_247;
  assign _T_3650 = release_state == 3'h7;
  assign _T_3651 = _T_3549 | _T_3650;
  assign _T_3653 = io_mem_0_c_bits_address[13:6];
  assign _T_3655 = metaArb_io_in_4_ready & metaArb_io_in_4_valid;
  assign _GEN_194 = _T_3655 ? 3'h0 : _GEN_192;
  assign _T_3657 = s1_valid | s2_valid;
  assign _T_3658 = _T_3657 | cached_grant_wait;
  assign _T_3661 = _T_3658 | uncachedInFlight_0;
  assign _T_3663 = _T_3661 == 1'h0;
  assign s1_xcpt_valid = tlb_io_req_valid & _T_146;
  assign _GEN_197 = s1_valid_not_nacked ? tlb_io_resp_pf_ld : _T_3669_pf_ld;
  assign _GEN_198 = s1_valid_not_nacked ? tlb_io_resp_pf_st : _T_3669_pf_st;
  assign _GEN_200 = s1_valid_not_nacked ? tlb_io_resp_ae_ld : _T_3669_ae_ld;
  assign _GEN_201 = s1_valid_not_nacked ? tlb_io_resp_ae_st : _T_3669_ae_st;
  assign _GEN_203 = s1_valid_not_nacked ? tlb_io_resp_ma_ld : _T_3669_ma_ld;
  assign _GEN_204 = s1_valid_not_nacked ? tlb_io_resp_ma_st : _T_3669_ma_st;
  assign _T_3687_pf_ld = _T_3667 ? _T_3669_pf_ld : 1'h0;
  assign _T_3687_pf_st = _T_3667 ? _T_3669_pf_st : 1'h0;
  assign _T_3687_ae_ld = _T_3667 ? _T_3669_ae_ld : 1'h0;
  assign _T_3687_ae_st = _T_3667 ? _T_3669_ae_st : 1'h0;
  assign _T_3687_ma_ld = _T_3667 ? _T_3669_ma_ld : 1'h0;
  assign _T_3687_ma_st = _T_3667 ? _T_3669_ma_st : 1'h0;
  assign _T_3690 = _T_3434 | s2_hit_valid;
  assign _T_3691 = _T_3690 | reset;
  assign _T_3693 = _T_3691 == 1'h0;
  assign _GEN_207 = s2_req_phys ? 1'h0 : _T_3687_ma_ld;
  assign _GEN_208 = s2_req_phys ? 1'h0 : _T_3687_ma_st;
  assign _GEN_209 = s2_req_phys ? 1'h0 : _T_3687_pf_ld;
  assign _GEN_210 = s2_req_phys ? 1'h0 : _T_3687_pf_st;
  assign _GEN_211 = s2_req_phys ? 1'h0 : _T_3687_ae_ld;
  assign _GEN_212 = s2_req_phys ? 1'h0 : _T_3687_ae_st;
  assign _T_3709 = _T_490 | _T_493;
  assign _T_3710 = s2_valid_masked & _T_3709;
  assign _T_3712 = _T_3710 == 1'h0;
  assign _T_3713 = _T_3712 | reset;
  assign _T_3715 = _T_3713 == 1'h0;
  assign _T_3717 = _T_3164 & _T_3197;
  assign _T_3721 = _T_1190 | reset;
  assign _T_3723 = _T_3721 == 1'h0;
  assign _GEN_213 = doUncachedResp ? 1'h1 : s2_valid_hit;
  assign _T_3726 = s2_req_typ[2];
  assign _T_3728 = _T_3726 == 1'h0;
  assign _T_3731 = s2_data_corrected[31:16];
  assign _T_3732 = s2_data_corrected[15:0];
  assign _T_3733 = _T_1809 ? _T_3731 : _T_3732;
  assign _T_3739 = _T_855 == 2'h1;
  assign _T_3741 = _T_3733[15];
  assign _T_3742 = _T_3728 & _T_3741;
  assign _T_3746 = _T_3742 ? 16'hffff : 16'h0;
  assign _T_3748 = _T_3739 ? _T_3746 : _T_3731;
  assign _T_3749 = {_T_3748,_T_3733};
  assign _T_3751 = _T_3749[15:8];
  assign _T_3752 = _T_3749[7:0];
  assign _T_3753 = _T_1819 ? _T_3751 : _T_3752;
  assign _T_3759 = _T_855 == 2'h0;
  assign _T_3761 = _T_3753[7];
  assign _T_3762 = _T_3728 & _T_3761;
  assign _T_3766 = _T_3762 ? 24'hffffff : 24'h0;
  assign _T_3767 = _T_3749[31:8];
  assign _T_3768 = _T_3759 ? _T_3766 : _T_3767;
  assign _T_3769 = {_T_3768,_T_3753};
  assign AMOALU_io_mask = pstore1_mask;
  assign AMOALU_io_cmd = pstore1_cmd;
  assign AMOALU_io_lhs = s2_data_corrected;
  assign AMOALU_io_rhs = a_data;
  assign _GEN_216 = AMOALU_io_out;
  assign flushCounterNext = flushCounter + 8'h1;
  assign _T_3780 = flushCounterNext[8:8];
  assign _T_3785 = _T_3158 & _T_900;
  assign _GEN_217 = _T_3785 ? 1'h0 : flushed;
  assign _T_3788 = s2_req_cmd == 5'h5;
  assign _T_3789 = s2_valid_masked & _T_3788;
  assign _T_3791 = flushed == 1'h0;
  assign _T_3800 = _T_898 & _T_905;
  assign _GEN_218 = _T_3791 ? _T_3800 : flushing;
  assign _GEN_219 = _T_3789 ? _T_3791 : _T_1201;
  assign _GEN_220 = _T_3789 ? _GEN_218 : flushing;
  assign _T_3801 = metaArb_io_in_5_ready & metaArb_io_in_5_valid;
  assign _T_3803 = s1_flush_valid == 1'h0;
  assign _T_3804 = _T_3801 & _T_3803;
  assign _T_3807 = _T_3804 & _T_910;
  assign _T_3809 = _T_3807 & _T_235;
  assign _T_3812 = _T_3809 & _T_898;
  assign _GEN_221 = _T_3780 ? 1'h1 : _GEN_217;
  assign _GEN_222 = s2_flush_valid_pre_tag_ecc ? flushCounterNext : {{1'd0}, flushCounter};
  assign _GEN_223 = s2_flush_valid_pre_tag_ecc ? _GEN_221 : _GEN_217;
  assign _T_3819 = flushed & _T_235;
  assign _T_3822 = _T_3819 & _T_898;
  assign _GEN_224 = _T_3822 ? 1'h0 : _GEN_220;
  assign _GEN_226 = flushing ? _GEN_222 : {{1'd0}, flushCounter};
  assign _GEN_227 = flushing ? _GEN_223 : _GEN_217;
  assign _GEN_228 = flushing ? _GEN_224 : _GEN_220;
  assign _GEN_229 = _T_3780 ? 1'h0 : resetting;
  assign _GEN_230 = resetting ? flushCounterNext : _GEN_226;
  assign _GEN_231 = resetting ? _GEN_229 : resetting;
  assign _GEN_248 = _T_3164 & grantIsCached;
  assign _GEN_250 = _T_3164 & _T_3230;
  assign _GEN_251 = _GEN_250 & _T_3238;
  assign _GEN_254 = _T_3164 & _T_3259;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  s1_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  s1_probe = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  probe_bits_param = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  probe_bits_address = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  s1_req_addr = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  s1_req_tag = _RAND_5[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  s1_req_cmd = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  s1_req_typ = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  s1_req_phys = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  s1_flush_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  cached_grant_wait = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  release_ack_wait = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  release_state = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  uncachedInFlight_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  uncachedReqs_0_addr = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  uncachedReqs_0_tag = _RAND_15[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  uncachedReqs_0_typ = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_461 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  s2_probe = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_478 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  s2_req_addr = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  s2_req_tag = _RAND_21[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  s2_req_cmd = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  s2_req_typ = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  s2_req_phys = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  s2_uncached = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  s2_flush_valid_pre_tag_ecc = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  s2_data = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  s2_probe_state_state = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  s2_hit_state_state = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  s2_waw_hazard = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_926_state = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  lrscCount = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  pstore1_cmd = _RAND_33[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  pstore1_addr = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  a_data = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  pstore1_mask = _RAND_36[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_1354 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  pstore2_valid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_1379 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  pstore2_addr = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_1422 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_1428 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_1434 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_1440 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  pstore2_storegen_mask = _RAND_45[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_3176 = _RAND_46[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  grantInProgress = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  blockProbeAfterGrantCount = _RAND_48[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  blockUncachedGrant = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_3454 = _RAND_50[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  s1_release_data_valid = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  s2_release_data_valid = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_3667 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_3669_pf_ld = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_3669_pf_st = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_3669_ae_ld = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_3669_ae_st = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_3669_ma_ld = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_3669_ma_st = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  doUncachedResp = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  resetting = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  flushed = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  flushing = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  flushCounter = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= _T_133;
    end
    if (reset) begin
      s1_probe <= 1'h0;
    end else begin
      if (_T_3539) begin
        if (metaArb_io_in_6_ready) begin
          s1_probe <= 1'h1;
        end else begin
          s1_probe <= _T_136;
        end
      end else begin
        s1_probe <= _T_136;
      end
    end
    if (_T_136) begin
      probe_bits_param <= io_mem_0_b_bits_param;
    end
    if (_T_136) begin
      probe_bits_address <= io_mem_0_b_bits_address;
    end
    if (_T_149) begin
      s1_req_addr <= _T_153;
    end
    if (_T_149) begin
      s1_req_tag <= io_cpu_req_bits_tag;
    end
    if (_T_149) begin
      s1_req_cmd <= io_cpu_req_bits_cmd;
    end
    if (_T_149) begin
      s1_req_typ <= io_cpu_req_bits_typ;
    end
    if (_T_149) begin
      s1_req_phys <= io_cpu_req_bits_phys;
    end
    s1_flush_valid <= _T_3812;
    if (reset) begin
      cached_grant_wait <= 1'h0;
    end else begin
      if (_T_3164) begin
        if (grantIsCached) begin
          if (d_last) begin
            cached_grant_wait <= 1'h0;
          end else begin
            if (_T_3158) begin
              if (_T_900) begin
                cached_grant_wait <= 1'h1;
              end
            end
          end
        end else begin
          if (_T_3158) begin
            if (_T_900) begin
              cached_grant_wait <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_3158) begin
          if (_T_900) begin
            cached_grant_wait <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      release_ack_wait <= 1'h0;
    end else begin
      if (_T_3550) begin
        if (_T_3636) begin
          release_ack_wait <= 1'h1;
        end else begin
          if (_T_3164) begin
            if (_T_3259) begin
              release_ack_wait <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_3164) begin
          if (_T_3259) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      release_state <= 3'h0;
    end else begin
      if (_T_3655) begin
        release_state <= 3'h0;
      end else begin
        if (_T_3550) begin
          if (_T_3441) begin
            release_state <= 3'h6;
          end else begin
            if (_T_233) begin
              if (_T_3441) begin
                release_state <= 3'h7;
              end else begin
                if (_T_3545) begin
                  if (_T_3441) begin
                    release_state <= 3'h7;
                  end else begin
                    if (_T_3543) begin
                      if (_T_3441) begin
                        release_state <= 3'h0;
                      end else begin
                        if (_T_3539) begin
                          if (metaArb_io_in_6_ready) begin
                            release_state <= 3'h0;
                          end else begin
                            if (s2_probe) begin
                              if (_T_3533) begin
                                if (_T_3441) begin
                                  release_state <= 3'h0;
                                end else begin
                                  release_state <= 3'h5;
                                end
                              end else begin
                                if (_T_3523) begin
                                  if (_T_3441) begin
                                    release_state <= 3'h7;
                                  end else begin
                                    release_state <= 3'h3;
                                  end
                                end else begin
                                  if (s2_prb_ack_data) begin
                                    release_state <= 3'h2;
                                  end
                                end
                              end
                            end
                          end
                        end else begin
                          if (s2_probe) begin
                            if (_T_3533) begin
                              if (_T_3441) begin
                                release_state <= 3'h0;
                              end else begin
                                release_state <= 3'h5;
                              end
                            end else begin
                              if (_T_3523) begin
                                if (_T_3441) begin
                                  release_state <= 3'h7;
                                end else begin
                                  release_state <= 3'h3;
                                end
                              end else begin
                                if (s2_prb_ack_data) begin
                                  release_state <= 3'h2;
                                end
                              end
                            end
                          end
                        end
                      end
                    end else begin
                      if (_T_3539) begin
                        if (metaArb_io_in_6_ready) begin
                          release_state <= 3'h0;
                        end else begin
                          if (s2_probe) begin
                            if (_T_3533) begin
                              if (_T_3441) begin
                                release_state <= 3'h0;
                              end else begin
                                release_state <= 3'h5;
                              end
                            end else begin
                              if (_T_3523) begin
                                if (_T_3441) begin
                                  release_state <= 3'h7;
                                end else begin
                                  release_state <= 3'h3;
                                end
                              end else begin
                                if (s2_prb_ack_data) begin
                                  release_state <= 3'h2;
                                end
                              end
                            end
                          end
                        end
                      end else begin
                        if (s2_probe) begin
                          if (_T_3533) begin
                            if (_T_3441) begin
                              release_state <= 3'h0;
                            end else begin
                              release_state <= 3'h5;
                            end
                          end else begin
                            if (_T_3523) begin
                              if (_T_3441) begin
                                release_state <= 3'h7;
                              end else begin
                                release_state <= 3'h3;
                              end
                            end else begin
                              if (s2_prb_ack_data) begin
                                release_state <= 3'h2;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_3543) begin
                    if (_T_3441) begin
                      release_state <= 3'h0;
                    end else begin
                      if (_T_3539) begin
                        if (metaArb_io_in_6_ready) begin
                          release_state <= 3'h0;
                        end else begin
                          release_state <= _GEN_143;
                        end
                      end else begin
                        release_state <= _GEN_143;
                      end
                    end
                  end else begin
                    if (_T_3539) begin
                      if (metaArb_io_in_6_ready) begin
                        release_state <= 3'h0;
                      end else begin
                        release_state <= _GEN_143;
                      end
                    end else begin
                      release_state <= _GEN_143;
                    end
                  end
                end
              end
            end else begin
              if (_T_3545) begin
                if (_T_3441) begin
                  release_state <= 3'h7;
                end else begin
                  if (_T_3543) begin
                    if (_T_3441) begin
                      release_state <= 3'h0;
                    end else begin
                      release_state <= _GEN_157;
                    end
                  end else begin
                    release_state <= _GEN_157;
                  end
                end
              end else begin
                if (_T_3543) begin
                  if (_T_3441) begin
                    release_state <= 3'h0;
                  end else begin
                    release_state <= _GEN_157;
                  end
                end else begin
                  release_state <= _GEN_157;
                end
              end
            end
          end
        end else begin
          if (_T_233) begin
            if (_T_3441) begin
              release_state <= 3'h7;
            end else begin
              if (_T_3545) begin
                if (_T_3441) begin
                  release_state <= 3'h7;
                end else begin
                  release_state <= _GEN_161;
                end
              end else begin
                release_state <= _GEN_161;
              end
            end
          end else begin
            if (_T_3545) begin
              if (_T_3441) begin
                release_state <= 3'h7;
              end else begin
                release_state <= _GEN_161;
              end
            end else begin
              release_state <= _GEN_161;
            end
          end
        end
      end
    end
    if (reset) begin
      uncachedInFlight_0 <= 1'h0;
    end else begin
      if (_T_3164) begin
        if (_T_3230) begin
          if (_T_3238) begin
            uncachedInFlight_0 <= 1'h0;
          end else begin
            if (_T_3158) begin
              if (s2_uncached) begin
                if (_T_3157) begin
                  uncachedInFlight_0 <= 1'h1;
                end
              end
            end
          end
        end else begin
          if (_T_3158) begin
            if (s2_uncached) begin
              if (_T_3157) begin
                uncachedInFlight_0 <= 1'h1;
              end
            end
          end
        end
      end else begin
        if (_T_3158) begin
          if (s2_uncached) begin
            if (_T_3157) begin
              uncachedInFlight_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (_T_3158) begin
      if (s2_uncached) begin
        if (_T_3157) begin
          uncachedReqs_0_addr <= s2_req_addr;
        end
      end
    end
    if (_T_3158) begin
      if (s2_uncached) begin
        if (_T_3157) begin
          uncachedReqs_0_tag <= s2_req_tag;
        end
      end
    end
    if (_T_3158) begin
      if (s2_uncached) begin
        if (_T_3157) begin
          uncachedReqs_0_typ <= s2_req_typ;
        end
      end
    end
    if (reset) begin
      _T_461 <= 1'h0;
    end else begin
      _T_461 <= _T_458;
    end
    if (reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    _T_478 <= _T_146;
    if (_T_3164) begin
      if (_T_3230) begin
        if (_T_3197) begin
          s2_req_addr <= _T_3253;
        end else begin
          if (_T_482) begin
            s2_req_addr <= tlb_io_resp_paddr;
          end
        end
      end else begin
        if (_T_482) begin
          s2_req_addr <= tlb_io_resp_paddr;
        end
      end
    end else begin
      if (_T_482) begin
        s2_req_addr <= tlb_io_resp_paddr;
      end
    end
    if (_T_3164) begin
      if (_T_3230) begin
        if (_T_3197) begin
          s2_req_tag <= uncachedReqs_0_tag;
        end else begin
          if (_T_482) begin
            s2_req_tag <= s1_req_tag;
          end
        end
      end else begin
        if (_T_482) begin
          s2_req_tag <= s1_req_tag;
        end
      end
    end else begin
      if (_T_482) begin
        s2_req_tag <= s1_req_tag;
      end
    end
    if (_T_3164) begin
      if (_T_3230) begin
        if (_T_3197) begin
          s2_req_cmd <= 5'h0;
        end else begin
          if (_T_482) begin
            s2_req_cmd <= s1_req_cmd;
          end
        end
      end else begin
        if (_T_482) begin
          s2_req_cmd <= s1_req_cmd;
        end
      end
    end else begin
      if (_T_482) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end
    if (_T_3164) begin
      if (_T_3230) begin
        if (_T_3197) begin
          s2_req_typ <= uncachedReqs_0_typ;
        end else begin
          if (_T_482) begin
            s2_req_typ <= s1_req_typ;
          end
        end
      end else begin
        if (_T_482) begin
          s2_req_typ <= s1_req_typ;
        end
      end
    end else begin
      if (_T_482) begin
        s2_req_typ <= s1_req_typ;
      end
    end
    if (_T_482) begin
      s2_req_phys <= s1_req_phys;
    end
    if (_T_482) begin
      s2_uncached <= 1'h1;
    end
    s2_flush_valid_pre_tag_ecc <= s1_flush_valid;
    if (_T_3164) begin
      if (_T_3230) begin
        if (_T_3197) begin
          s2_data <= _T_3249;
        end else begin
          if (_T_571) begin
            s2_data <= data_io_resp_0;
          end
        end
      end else begin
        if (_T_571) begin
          s2_data <= data_io_resp_0;
        end
      end
    end else begin
      if (_T_571) begin
        s2_data <= data_io_resp_0;
      end
    end
    if (s1_probe) begin
      if (s1_hit_way) begin
        s2_probe_state_state <= 2'h3;
      end else begin
        s2_probe_state_state <= 2'h0;
      end
    end
    if (s1_valid_not_nacked) begin
      if (s1_hit_way) begin
        s2_hit_state_state <= 2'h3;
      end else begin
        s2_hit_state_state <= 2'h0;
      end
    end
    if (s1_valid_not_nacked) begin
      s2_waw_hazard <= 1'h0;
    end
    if (_T_482) begin
      _T_926_state <= 2'h0;
    end
    if (reset) begin
      lrscCount <= 5'h0;
    end else begin
      if (_T_1256) begin
        lrscCount <= 5'h0;
      end else begin
        if (_T_1248) begin
          lrscCount <= _T_1252;
        end
      end
    end
    if (_T_1262) begin
      pstore1_cmd <= s1_req_cmd;
    end
    if (_T_1262) begin
      pstore1_addr <= tlb_io_resp_paddr;
    end
    if (_T_1262) begin
      a_data <= io_cpu_s1_data_data;
    end
    if (_T_1262) begin
      if (_T_191) begin
        pstore1_mask <= io_cpu_s1_data_mask;
      end else begin
        pstore1_mask <= _T_455;
      end
    end
    if (_T_1262) begin
      _T_1354 <= _T_1351;
    end
    pstore2_valid <= _T_1402;
    _T_1379 <= _T_1395;
    if (advance_pstore1) begin
      pstore2_addr <= pstore1_addr;
    end
    if (advance_pstore1) begin
      _T_1422 <= _T_1417;
    end
    if (advance_pstore1) begin
      _T_1428 <= _T_1423;
    end
    if (advance_pstore1) begin
      _T_1434 <= _T_1429;
    end
    if (advance_pstore1) begin
      _T_1440 <= _T_1435;
    end
    if (advance_pstore1) begin
      pstore2_storegen_mask <= _T_1451;
    end
    if (reset) begin
      _T_3176 <= 10'h0;
    end else begin
      if (_T_3164) begin
        if (d_first) begin
          if (_T_3171) begin
            _T_3176 <= _T_3170;
          end else begin
            _T_3176 <= 10'h0;
          end
        end else begin
          _T_3176 <= _T_3180;
        end
      end
    end
    if (reset) begin
      grantInProgress <= 1'h0;
    end else begin
      if (_T_3164) begin
        if (grantIsCached) begin
          if (d_last) begin
            grantInProgress <= 1'h0;
          end else begin
            grantInProgress <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      blockProbeAfterGrantCount <= 3'h0;
    end else begin
      if (_T_3164) begin
        if (grantIsCached) begin
          if (d_last) begin
            blockProbeAfterGrantCount <= 3'h7;
          end else begin
            if (_T_3208) begin
              blockProbeAfterGrantCount <= _T_3212;
            end
          end
        end else begin
          if (_T_3208) begin
            blockProbeAfterGrantCount <= _T_3212;
          end
        end
      end else begin
        if (_T_3208) begin
          blockProbeAfterGrantCount <= _T_3212;
        end
      end
    end
    if (_T_3401) begin
      if (io_mem_0_d_valid) begin
        blockUncachedGrant <= _T_3267;
      end else begin
        blockUncachedGrant <= dataArb_io_out_valid;
      end
    end else begin
      blockUncachedGrant <= dataArb_io_out_valid;
    end
    if (reset) begin
      _T_3454 <= 10'h0;
    end else begin
      if (_T_3441) begin
        if (c_first) begin
          _T_3454 <= 10'h0;
        end else begin
          _T_3454 <= _T_3458;
        end
      end
    end
    s1_release_data_valid <= _T_3468;
    s2_release_data_valid <= _T_3472;
    _T_3667 <= s1_xcpt_valid;
    if (s1_valid_not_nacked) begin
      _T_3669_pf_ld <= tlb_io_resp_pf_ld;
    end
    if (s1_valid_not_nacked) begin
      _T_3669_pf_st <= tlb_io_resp_pf_st;
    end
    if (s1_valid_not_nacked) begin
      _T_3669_ae_ld <= tlb_io_resp_ae_ld;
    end
    if (s1_valid_not_nacked) begin
      _T_3669_ae_st <= tlb_io_resp_ae_st;
    end
    if (s1_valid_not_nacked) begin
      _T_3669_ma_ld <= tlb_io_resp_ma_ld;
    end
    if (s1_valid_not_nacked) begin
      _T_3669_ma_st <= tlb_io_resp_ma_st;
    end
    doUncachedResp <= io_cpu_replay_next;
    if (reset) begin
      resetting <= 1'h1;
    end else begin
      if (resetting) begin
        if (_T_3780) begin
          resetting <= 1'h0;
        end
      end
    end
    if (reset) begin
      flushed <= 1'h1;
    end else begin
      if (flushing) begin
        if (s2_flush_valid_pre_tag_ecc) begin
          if (_T_3780) begin
            flushed <= 1'h1;
          end else begin
            if (_T_3785) begin
              flushed <= 1'h0;
            end
          end
        end else begin
          if (_T_3785) begin
            flushed <= 1'h0;
          end
        end
      end else begin
        if (_T_3785) begin
          flushed <= 1'h0;
        end
      end
    end
    if (reset) begin
      flushing <= 1'h0;
    end else begin
      if (flushing) begin
        if (_T_3822) begin
          flushing <= 1'h0;
        end else begin
          if (_T_3789) begin
            if (_T_3791) begin
              flushing <= _T_3800;
            end
          end
        end
      end else begin
        if (_T_3789) begin
          if (_T_3791) begin
            flushing <= _T_3800;
          end
        end
      end
    end
    if (reset) begin
      flushCounter <= 8'h0;
    end else begin
      flushCounter <= _GEN_230[7:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1387) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:296 assert(!s2_store_valid || !pstore1_held)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_248 & _T_3223) begin
          $fwrite(32'h80000002,"Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:404 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_248 & _T_3223) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_251 & _T_3241) begin
          $fwrite(32'h80000002,"Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:416 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_251 & _T_3241) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_254 & _T_3262) begin
          $fwrite(32'h80000002,"Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:429 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_254 & _T_3262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3282) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:447 assert(!metaArb.io.in(3).valid || metaArb.io.in(3).ready)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3282) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3413 & _T_3417) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:470 when (tl_out.e.fire()) { assert(tl_out.d.fire()) }\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3413 & _T_3417) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:498 assert(!(s2_valid && s2_hit_valid && !s2_data_error))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_req_phys & _T_3693) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:584 assert(!s2_valid || s2_hit_valid)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (s2_req_phys & _T_3693) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3715) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:587 assert(!(s2_valid_masked && s2_req.cmd.isOneOf(M_XLR, M_XSC)))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_3715) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & _T_3723) begin
          $fwrite(32'h80000002,"Assertion failed\n    at DCache.scala:594 assert(!s2_valid_hit)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & _T_3723) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ICache_icache(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [31:0] io_req_bits_addr,
  input  [31:0] io_s1_paddr,
  input         io_s1_kill,
  input         io_s2_kill,
  output        io_resp_valid,
  output [31:0] io_resp_bits_data,
  output        io_resp_bits_ae,
  input         io_invalidate,
  input         io_tl_out_0_a_ready,
  output        io_tl_out_0_a_valid,
  output [2:0]  io_tl_out_0_a_bits_opcode,
  output [2:0]  io_tl_out_0_a_bits_param,
  output [3:0]  io_tl_out_0_a_bits_size,
  output        io_tl_out_0_a_bits_source,
  output [31:0] io_tl_out_0_a_bits_address,
  output [3:0]  io_tl_out_0_a_bits_mask,
  output [31:0] io_tl_out_0_a_bits_data,
  output        io_tl_out_0_d_ready,
  input         io_tl_out_0_d_valid,
  input  [2:0]  io_tl_out_0_d_bits_opcode,
  input  [3:0]  io_tl_out_0_d_bits_size,
  input  [31:0] io_tl_out_0_d_bits_data,
  input         io_tl_out_0_d_bits_error
);
  reg  s1_slaveValid;
  reg [31:0] _RAND_0;
  reg  s3_slaveValid;
  reg [31:0] _RAND_1;
  reg  s1_valid;
  reg [31:0] _RAND_2;
  wire  s1_hit;
  wire  _T_67;
  wire  _T_68;
  reg  s2_valid;
  reg [31:0] _RAND_3;
  reg  s2_hit;
  reg [31:0] _RAND_4;
  reg  invalidated;
  reg [31:0] _RAND_5;
  reg  refill_valid;
  reg [31:0] _RAND_6;
  wire  _T_76;
  wire  _T_77;
  wire  _T_79;
  wire  _T_80;
  reg  _T_82;
  reg [31:0] _RAND_7;
  wire  _T_84;
  wire  s2_miss;
  wire  _T_85;
  wire  _T_87;
  wire  _T_88;
  reg [31:0] refill_addr;
  reg [31:0] _RAND_8;
  wire [31:0] _GEN_0;
  wire [19:0] refill_tag;
  wire [5:0] refill_idx;
  wire  _T_90;
  wire  _T_92;
  wire  _T_94;
  wire  s0_valid;
  wire [26:0] _T_98;
  wire [11:0] _T_99;
  wire [11:0] _T_100;
  wire [9:0] _T_101;
  wire  _T_102;
  wire [9:0] _T_104;
  reg [9:0] _T_107;
  reg [31:0] _RAND_9;
  wire [10:0] _T_109;
  wire [10:0] _T_110;
  wire [9:0] _T_111;
  wire  _T_113;
  wire  _T_115;
  wire  _T_117;
  wire  _T_118;
  wire  refill_done;
  wire [9:0] _T_119;
  wire [9:0] refill_cnt;
  wire [9:0] _T_120;
  wire [9:0] _GEN_1;
  wire  _T_122;
  wire [5:0] tag_array_RW0_addr;
  wire  tag_array_RW0_en;
  wire  tag_array_RW0_clk;
  wire  tag_array_RW0_wmode;
  wire [20:0] tag_array_RW0_wdata_0;
  wire [20:0] tag_array_RW0_rdata_0;
  wire  tag_array_RW0_wmask_0;
  wire [5:0] _T_130;
  wire  _T_132;
  wire  _T_133;
  reg  accruedRefillError;
  reg [31:0] _RAND_10;
  wire  _T_146;
  wire  _T_147;
  wire  refillError;
  wire [20:0] _T_148;
  reg [63:0] vb_array;
  reg [63:0] _RAND_11;
  wire [6:0] _T_166;
  wire  _T_168;
  wire  _T_169;
  wire [127:0] _T_171;
  wire [127:0] _GEN_37;
  wire [127:0] _T_172;
  wire [63:0] _T_173;
  wire [127:0] _GEN_38;
  wire [127:0] _T_174;
  wire [127:0] _T_175;
  wire [127:0] _T_176;
  wire  _GEN_13;
  wire [127:0] _GEN_14;
  wire [127:0] _GEN_15;
  wire  _GEN_16;
  reg [11:0] s1s3_slaveAddr;
  reg [31:0] _RAND_12;
  reg [31:0] s1s3_slaveData;
  reg [31:0] _RAND_13;
  wire [5:0] _T_200;
  wire [19:0] _T_201;
  wire [6:0] _T_222;
  wire [63:0] _T_223;
  wire  _T_224;
  wire  _T_226;
  wire  _T_227;
  wire  _T_228;
  wire [19:0] _T_229;
  wire  _T_230;
  wire  _T_231;
  wire  _T_237;
  wire  _T_239;
  wire [9:0] data_arrays_0_RW0_addr;
  wire  data_arrays_0_RW0_en;
  wire  data_arrays_0_RW0_clk;
  wire  data_arrays_0_RW0_wmode;
  wire [31:0] data_arrays_0_RW0_wdata_0;
  wire [31:0] data_arrays_0_RW0_rdata_0;
  wire  data_arrays_0_RW0_wmask_0;
  wire  _T_270;
  wire  _T_275;
  wire [9:0] _GEN_39;
  wire [9:0] _T_277;
  wire [9:0] _T_278;
  wire [9:0] _T_279;
  wire [9:0] _T_281;
  wire [9:0] _T_283;
  wire [9:0] _T_284;
  wire [31:0] _T_286;
  wire  _T_304;
  wire  _T_305;
  wire [31:0] _GEN_28;
  reg [31:0] _T_343_0;
  reg [31:0] _RAND_14;
  wire [31:0] _GEN_30;
  reg  _T_358_0;
  reg [31:0] _RAND_15;
  wire  _GEN_31;
  reg  _T_372;
  reg [31:0] _RAND_16;
  wire  _GEN_32;
  wire  _T_377;
  wire  _GEN_33;
  wire  _T_379;
  wire  _T_381;
  wire  _T_382;
  wire  _T_384;
  wire  _T_385;
  wire [25:0] _T_387;
  wire [31:0] _GEN_40;
  wire [31:0] _T_388;
  wire  _GEN_34;
  wire  _T_526;
  wire  _GEN_35;
  wire  _GEN_36;
  tag_array tag_array (
    .RW0_addr(tag_array_RW0_addr),
    .RW0_en(tag_array_RW0_en),
    .RW0_clk(tag_array_RW0_clk),
    .RW0_wmode(tag_array_RW0_wmode),
    .RW0_wdata_0(tag_array_RW0_wdata_0),
    .RW0_rdata_0(tag_array_RW0_rdata_0),
    .RW0_wmask_0(tag_array_RW0_wmask_0)
  );
  data_arrays_0_0 data_arrays_0 (
    .RW0_addr(data_arrays_0_RW0_addr),
    .RW0_en(data_arrays_0_RW0_en),
    .RW0_clk(data_arrays_0_RW0_clk),
    .RW0_wmode(data_arrays_0_RW0_wmode),
    .RW0_wdata_0(data_arrays_0_RW0_wdata_0),
    .RW0_rdata_0(data_arrays_0_RW0_rdata_0),
    .RW0_wmask_0(data_arrays_0_RW0_wmask_0)
  );
  assign io_req_ready = _T_94;
  assign io_resp_valid = _T_382;
  assign io_resp_bits_data = _T_343_0;
  assign io_resp_bits_ae = _T_372;
  assign io_tl_out_0_a_valid = _T_385;
  assign io_tl_out_0_a_bits_opcode = 3'h4;
  assign io_tl_out_0_a_bits_param = 3'h0;
  assign io_tl_out_0_a_bits_size = 4'h6;
  assign io_tl_out_0_a_bits_source = 1'h0;
  assign io_tl_out_0_a_bits_address = _T_388;
  assign io_tl_out_0_a_bits_mask = 4'hf;
  assign io_tl_out_0_a_bits_data = 32'h0;
  assign io_tl_out_0_d_ready = _T_122;
  assign s1_hit = _T_231 | s1_slaveValid;
  assign _T_67 = io_s1_kill == 1'h0;
  assign _T_68 = s1_valid & _T_67;
  assign _T_76 = s2_hit == 1'h0;
  assign _T_77 = s2_valid & _T_76;
  assign _T_79 = io_s2_kill == 1'h0;
  assign _T_80 = _T_77 & _T_79;
  assign _T_84 = _T_82 == 1'h0;
  assign s2_miss = _T_80 & _T_84;
  assign _T_85 = refill_valid | s2_miss;
  assign _T_87 = _T_85 == 1'h0;
  assign _T_88 = s1_valid & _T_87;
  assign _GEN_0 = _T_88 ? io_s1_paddr : refill_addr;
  assign refill_tag = refill_addr[31:12];
  assign refill_idx = refill_addr[11:6];
  assign _T_90 = io_tl_out_0_d_ready & io_tl_out_0_d_valid;
  assign _T_92 = _T_90 | s3_slaveValid;
  assign _T_94 = _T_92 == 1'h0;
  assign s0_valid = io_req_ready & io_req_valid;
  assign _T_98 = 27'hfff << io_tl_out_0_d_bits_size;
  assign _T_99 = _T_98[11:0];
  assign _T_100 = ~ _T_99;
  assign _T_101 = _T_100[11:2];
  assign _T_102 = io_tl_out_0_d_bits_opcode[0];
  assign _T_104 = _T_102 ? _T_101 : 10'h0;
  assign _T_109 = _T_107 - 10'h1;
  assign _T_110 = $unsigned(_T_109);
  assign _T_111 = _T_110[9:0];
  assign _T_113 = _T_107 == 10'h0;
  assign _T_115 = _T_107 == 10'h1;
  assign _T_117 = _T_104 == 10'h0;
  assign _T_118 = _T_115 | _T_117;
  assign refill_done = _T_118 & _T_90;
  assign _T_119 = ~ _T_111;
  assign refill_cnt = _T_104 & _T_119;
  assign _T_120 = _T_113 ? _T_104 : _T_111;
  assign _GEN_1 = _T_90 ? _T_120 : _T_107;
  assign _T_122 = s3_slaveValid == 1'h0;
  assign tag_array_RW0_addr = refill_done ? refill_idx : _T_130;
  assign tag_array_RW0_en = _T_133 | refill_done;
  assign tag_array_RW0_clk = clock;
  assign tag_array_RW0_wmode = refill_done;
  assign tag_array_RW0_wdata_0 = _T_148;
  assign tag_array_RW0_wmask_0 = refill_done;
  assign _T_130 = io_req_bits_addr[11:6];
  assign _T_132 = refill_done == 1'h0;
  assign _T_133 = _T_132 & s0_valid;
  assign _T_146 = refill_cnt > 10'h0;
  assign _T_147 = _T_146 & accruedRefillError;
  assign refillError = io_tl_out_0_d_bits_error | _T_147;
  assign _T_148 = {refillError,refill_tag};
  assign _T_166 = {1'h0,refill_idx};
  assign _T_168 = invalidated == 1'h0;
  assign _T_169 = refill_done & _T_168;
  assign _T_171 = 128'h1 << _T_166;
  assign _GEN_37 = {{64'd0}, vb_array};
  assign _T_172 = _GEN_37 | _T_171;
  assign _T_173 = ~ vb_array;
  assign _GEN_38 = {{64'd0}, _T_173};
  assign _T_174 = _GEN_38 | _T_171;
  assign _T_175 = ~ _T_174;
  assign _T_176 = _T_169 ? _T_172 : _T_175;
  assign _GEN_13 = _T_90 ? refillError : accruedRefillError;
  assign _GEN_14 = _T_90 ? _T_176 : {{64'd0}, vb_array};
  assign _GEN_15 = _GEN_33 ? 128'h0 : _GEN_14;
  assign _GEN_16 = _GEN_33 ? 1'h1 : invalidated;
  assign _T_200 = io_s1_paddr[11:6];
  assign _T_201 = io_s1_paddr[31:12];
  assign _T_222 = {1'h0,_T_200};
  assign _T_223 = vb_array >> _T_222;
  assign _T_224 = _T_223[0];
  assign _T_226 = s1_slaveValid == 1'h0;
  assign _T_227 = _T_224 & _T_226;
  assign _T_228 = tag_array_RW0_rdata_0[20];
  assign _T_229 = tag_array_RW0_rdata_0[19:0];
  assign _T_230 = _T_229 == _T_201;
  assign _T_231 = _T_227 & _T_230;
  assign _T_237 = _T_231 & _T_228;
  assign _T_239 = s1_valid | s1_slaveValid;
  assign data_arrays_0_RW0_addr = _T_284;
  assign data_arrays_0_RW0_en = _T_305 | _T_275;
  assign data_arrays_0_RW0_clk = clock;
  assign data_arrays_0_RW0_wmode = _T_275;
  assign data_arrays_0_RW0_wdata_0 = _T_286;
  assign data_arrays_0_RW0_wmask_0 = _T_275;
  assign _T_270 = _T_90 & _T_168;
  assign _T_275 = _T_270 | s3_slaveValid;
  assign _GEN_39 = {{4'd0}, refill_idx};
  assign _T_277 = _GEN_39 << 4;
  assign _T_278 = _T_277 | refill_cnt;
  assign _T_279 = s1s3_slaveAddr[11:2];
  assign _T_281 = io_req_bits_addr[11:2];
  assign _T_283 = s3_slaveValid ? _T_279 : _T_281;
  assign _T_284 = _T_90 ? _T_278 : _T_283;
  assign _T_286 = s3_slaveValid ? s1s3_slaveData : io_tl_out_0_d_bits_data;
  assign _T_304 = _T_275 == 1'h0;
  assign _T_305 = _T_304 & s0_valid;
  assign _GEN_28 = data_arrays_0_RW0_rdata_0;
  assign _GEN_30 = _T_239 ? _GEN_28 : _T_343_0;
  assign _GEN_31 = _T_239 ? 1'h0 : _T_358_0;
  assign _GEN_32 = _T_239 ? _T_237 : _T_372;
  assign _T_377 = s2_valid & _T_358_0;
  assign _GEN_33 = _T_377 ? 1'h1 : io_invalidate;
  assign _T_379 = s2_valid & s2_hit;
  assign _T_381 = _T_358_0 == 1'h0;
  assign _T_382 = _T_379 & _T_381;
  assign _T_384 = refill_valid == 1'h0;
  assign _T_385 = s2_miss & _T_384;
  assign _T_387 = refill_addr[31:6];
  assign _GEN_40 = {{6'd0}, _T_387};
  assign _T_388 = _GEN_40 << 6;
  assign _GEN_34 = _T_384 ? 1'h0 : _GEN_16;
  assign _T_526 = io_tl_out_0_a_ready & io_tl_out_0_a_valid;
  assign _GEN_35 = _T_526 ? 1'h1 : refill_valid;
  assign _GEN_36 = refill_done ? 1'h0 : _GEN_35;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  s1_slaveValid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  s3_slaveValid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  s1_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  s2_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  s2_hit = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  invalidated = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  refill_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_82 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  refill_addr = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_107 = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  accruedRefillError = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{$random}};
  vb_array = _RAND_11[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  s1s3_slaveAddr = _RAND_12[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  s1s3_slaveData = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_343_0 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_358_0 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_372 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      s1_slaveValid <= 1'h0;
    end else begin
      s1_slaveValid <= 1'h0;
    end
    s3_slaveValid <= 1'h0;
    if (reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= s0_valid;
    end
    if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _T_68;
    end
    s2_hit <= s1_hit;
    if (_T_384) begin
      invalidated <= 1'h0;
    end else begin
      if (_GEN_33) begin
        invalidated <= 1'h1;
      end
    end
    if (reset) begin
      refill_valid <= 1'h0;
    end else begin
      if (refill_done) begin
        refill_valid <= 1'h0;
      end else begin
        if (_T_526) begin
          refill_valid <= 1'h1;
        end
      end
    end
    _T_82 <= refill_valid;
    if (_T_88) begin
      refill_addr <= io_s1_paddr;
    end
    if (reset) begin
      _T_107 <= 10'h0;
    end else begin
      if (_T_90) begin
        if (_T_113) begin
          if (_T_102) begin
            _T_107 <= _T_101;
          end else begin
            _T_107 <= 10'h0;
          end
        end else begin
          _T_107 <= _T_111;
        end
      end
    end
    if (_T_90) begin
      accruedRefillError <= refillError;
    end
    if (reset) begin
      vb_array <= 64'h0;
    end else begin
      vb_array <= _GEN_15[63:0];
    end
    if (_T_239) begin
      _T_343_0 <= _GEN_28;
    end
    if (_T_239) begin
      _T_358_0 <= 1'h0;
    end
    if (_T_239) begin
      _T_372 <= _T_237;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ICache.scala:200 assert(!(s1_valid || s1_slaveValid) || PopCount(s1_tag_hit zip s1_tag_disparity map { case (h, d) => h && !d }) <= 1)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ICache.scala:306 assert(!(tl_out.a.valid && addrMaybeInScratchpad(tl_out.a.bits.address)))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ShiftQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_btb_valid,
  input         io_enq_bits_btb_bits_taken,
  input         io_enq_bits_btb_bits_bridx,
  input  [31:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_xcpt_pf_inst,
  input         io_enq_bits_xcpt_ae_inst,
  input         io_enq_bits_replay,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_btb_valid,
  output        io_deq_bits_btb_bits_taken,
  output        io_deq_bits_btb_bits_bridx,
  output [31:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_xcpt_pf_inst,
  output        io_deq_bits_xcpt_ae_inst,
  output        io_deq_bits_replay,
  output [4:0]  io_mask
);
  reg  valid_0;
  reg [31:0] _RAND_0;
  reg  valid_1;
  reg [31:0] _RAND_1;
  reg  valid_2;
  reg [31:0] _RAND_2;
  reg  valid_3;
  reg [31:0] _RAND_3;
  reg  valid_4;
  reg [31:0] _RAND_4;
  reg  elts_0_btb_valid;
  reg [31:0] _RAND_5;
  reg  elts_0_btb_bits_taken;
  reg [31:0] _RAND_6;
  reg  elts_0_btb_bits_bridx;
  reg [31:0] _RAND_7;
  reg [31:0] elts_0_pc;
  reg [31:0] _RAND_8;
  reg [31:0] elts_0_data;
  reg [31:0] _RAND_9;
  reg  elts_0_xcpt_pf_inst;
  reg [31:0] _RAND_10;
  reg  elts_0_xcpt_ae_inst;
  reg [31:0] _RAND_11;
  reg  elts_0_replay;
  reg [31:0] _RAND_12;
  reg  elts_1_btb_valid;
  reg [31:0] _RAND_13;
  reg  elts_1_btb_bits_taken;
  reg [31:0] _RAND_14;
  reg  elts_1_btb_bits_bridx;
  reg [31:0] _RAND_15;
  reg [31:0] elts_1_pc;
  reg [31:0] _RAND_16;
  reg [31:0] elts_1_data;
  reg [31:0] _RAND_17;
  reg  elts_1_xcpt_pf_inst;
  reg [31:0] _RAND_18;
  reg  elts_1_xcpt_ae_inst;
  reg [31:0] _RAND_19;
  reg  elts_1_replay;
  reg [31:0] _RAND_20;
  reg  elts_2_btb_valid;
  reg [31:0] _RAND_21;
  reg  elts_2_btb_bits_taken;
  reg [31:0] _RAND_22;
  reg  elts_2_btb_bits_bridx;
  reg [31:0] _RAND_23;
  reg [31:0] elts_2_pc;
  reg [31:0] _RAND_24;
  reg [31:0] elts_2_data;
  reg [31:0] _RAND_25;
  reg  elts_2_xcpt_pf_inst;
  reg [31:0] _RAND_26;
  reg  elts_2_xcpt_ae_inst;
  reg [31:0] _RAND_27;
  reg  elts_2_replay;
  reg [31:0] _RAND_28;
  reg  elts_3_btb_valid;
  reg [31:0] _RAND_29;
  reg  elts_3_btb_bits_taken;
  reg [31:0] _RAND_30;
  reg  elts_3_btb_bits_bridx;
  reg [31:0] _RAND_31;
  reg [31:0] elts_3_pc;
  reg [31:0] _RAND_32;
  reg [31:0] elts_3_data;
  reg [31:0] _RAND_33;
  reg  elts_3_xcpt_pf_inst;
  reg [31:0] _RAND_34;
  reg  elts_3_xcpt_ae_inst;
  reg [31:0] _RAND_35;
  reg  elts_3_replay;
  reg [31:0] _RAND_36;
  reg  elts_4_btb_valid;
  reg [31:0] _RAND_37;
  reg  elts_4_btb_bits_taken;
  reg [31:0] _RAND_38;
  reg  elts_4_btb_bits_bridx;
  reg [31:0] _RAND_39;
  reg [31:0] elts_4_pc;
  reg [31:0] _RAND_40;
  reg [31:0] elts_4_data;
  reg [31:0] _RAND_41;
  reg  elts_4_xcpt_pf_inst;
  reg [31:0] _RAND_42;
  reg  elts_4_xcpt_ae_inst;
  reg [31:0] _RAND_43;
  reg  elts_4_replay;
  reg [31:0] _RAND_44;
  wire  do_enq;
  wire  do_deq;
  wire  _T_143_btb_valid;
  wire  _T_143_btb_bits_taken;
  wire  _T_143_btb_bits_bridx;
  wire [31:0] _T_143_pc;
  wire [31:0] _T_143_data;
  wire  _T_143_xcpt_pf_inst;
  wire  _T_143_xcpt_ae_inst;
  wire  _T_143_replay;
  wire  _T_147;
  wire  _T_150;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire  _GEN_0;
  wire  _GEN_2;
  wire  _GEN_4;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _T_156_btb_valid;
  wire  _T_156_btb_bits_taken;
  wire  _T_156_btb_bits_bridx;
  wire [31:0] _T_156_pc;
  wire [31:0] _T_156_data;
  wire  _T_156_xcpt_pf_inst;
  wire  _T_156_xcpt_ae_inst;
  wire  _T_156_replay;
  wire  _T_160;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _T_166;
  wire  _T_167;
  wire  _GEN_16;
  wire  _GEN_18;
  wire  _GEN_20;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _T_168_btb_valid;
  wire  _T_168_btb_bits_taken;
  wire  _T_168_btb_bits_bridx;
  wire [31:0] _T_168_pc;
  wire [31:0] _T_168_data;
  wire  _T_168_xcpt_pf_inst;
  wire  _T_168_xcpt_ae_inst;
  wire  _T_168_replay;
  wire  _T_172;
  wire  _T_175;
  wire  _T_176;
  wire  _T_177;
  wire  _T_178;
  wire  _T_179;
  wire  _GEN_32;
  wire  _GEN_34;
  wire  _GEN_36;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _T_180_btb_valid;
  wire  _T_180_btb_bits_taken;
  wire  _T_180_btb_bits_bridx;
  wire [31:0] _T_180_pc;
  wire [31:0] _T_180_data;
  wire  _T_180_xcpt_pf_inst;
  wire  _T_180_xcpt_ae_inst;
  wire  _T_180_replay;
  wire  _T_184;
  wire  _T_187;
  wire  _T_188;
  wire  _T_189;
  wire  _T_190;
  wire  _T_191;
  wire  _GEN_48;
  wire  _GEN_50;
  wire  _GEN_52;
  wire [31:0] _GEN_58;
  wire [31:0] _GEN_59;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _T_195;
  wire  _T_196;
  wire  _T_197;
  wire  _T_198;
  wire  _GEN_64;
  wire  _GEN_66;
  wire  _GEN_68;
  wire [31:0] _GEN_74;
  wire [31:0] _GEN_75;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _T_201;
  wire  _T_202;
  wire  _GEN_80;
  wire  _T_206;
  wire  _T_207;
  wire  _T_210;
  wire  _GEN_81;
  wire  _T_215;
  wire  _GEN_82;
  wire  _T_222;
  wire  _GEN_83;
  wire  _T_227;
  wire  _GEN_84;
  wire  _T_234;
  wire  _GEN_85;
  wire  _T_239;
  wire  _GEN_86;
  wire  _T_246;
  wire  _GEN_87;
  wire  _T_251;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _GEN_91;
  wire  _GEN_93;
  wire  _GEN_95;
  wire [31:0] _GEN_101;
  wire [31:0] _GEN_102;
  wire  _GEN_104;
  wire  _GEN_105;
  wire  _GEN_106;
  wire [1:0] _T_265;
  wire [1:0] _T_266;
  wire [2:0] _T_267;
  wire [4:0] _T_268;
  assign io_enq_ready = _T_195;
  assign io_deq_valid = _GEN_90;
  assign io_deq_bits_btb_valid = _GEN_91;
  assign io_deq_bits_btb_bits_taken = _GEN_93;
  assign io_deq_bits_btb_bits_bridx = _GEN_95;
  assign io_deq_bits_pc = _GEN_101;
  assign io_deq_bits_data = _GEN_102;
  assign io_deq_bits_xcpt_pf_inst = _GEN_104;
  assign io_deq_bits_xcpt_ae_inst = _GEN_105;
  assign io_deq_bits_replay = _GEN_106;
  assign io_mask = _T_268;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign _T_143_btb_valid = valid_1 ? elts_1_btb_valid : io_enq_bits_btb_valid;
  assign _T_143_btb_bits_taken = valid_1 ? elts_1_btb_bits_taken : io_enq_bits_btb_bits_taken;
  assign _T_143_btb_bits_bridx = valid_1 ? elts_1_btb_bits_bridx : io_enq_bits_btb_bits_bridx;
  assign _T_143_pc = valid_1 ? elts_1_pc : io_enq_bits_pc;
  assign _T_143_data = valid_1 ? elts_1_data : io_enq_bits_data;
  assign _T_143_xcpt_pf_inst = valid_1 ? elts_1_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst;
  assign _T_143_xcpt_ae_inst = valid_1 ? elts_1_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst;
  assign _T_143_replay = valid_1 ? elts_1_replay : io_enq_bits_replay;
  assign _T_147 = io_deq_ready & valid_1;
  assign _T_150 = valid_0 == 1'h0;
  assign _T_153 = io_deq_ready ? valid_0 : _T_150;
  assign _T_154 = do_enq & _T_153;
  assign _T_155 = _T_147 | _T_154;
  assign _GEN_0 = _T_155 ? _T_143_btb_valid : elts_0_btb_valid;
  assign _GEN_2 = _T_155 ? _T_143_btb_bits_taken : elts_0_btb_bits_taken;
  assign _GEN_4 = _T_155 ? _T_143_btb_bits_bridx : elts_0_btb_bits_bridx;
  assign _GEN_10 = _T_155 ? _T_143_pc : elts_0_pc;
  assign _GEN_11 = _T_155 ? _T_143_data : elts_0_data;
  assign _GEN_13 = _T_155 ? _T_143_xcpt_pf_inst : elts_0_xcpt_pf_inst;
  assign _GEN_14 = _T_155 ? _T_143_xcpt_ae_inst : elts_0_xcpt_ae_inst;
  assign _GEN_15 = _T_155 ? _T_143_replay : elts_0_replay;
  assign _T_156_btb_valid = valid_2 ? elts_2_btb_valid : io_enq_bits_btb_valid;
  assign _T_156_btb_bits_taken = valid_2 ? elts_2_btb_bits_taken : io_enq_bits_btb_bits_taken;
  assign _T_156_btb_bits_bridx = valid_2 ? elts_2_btb_bits_bridx : io_enq_bits_btb_bits_bridx;
  assign _T_156_pc = valid_2 ? elts_2_pc : io_enq_bits_pc;
  assign _T_156_data = valid_2 ? elts_2_data : io_enq_bits_data;
  assign _T_156_xcpt_pf_inst = valid_2 ? elts_2_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst;
  assign _T_156_xcpt_ae_inst = valid_2 ? elts_2_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst;
  assign _T_156_replay = valid_2 ? elts_2_replay : io_enq_bits_replay;
  assign _T_160 = io_deq_ready & valid_2;
  assign _T_163 = valid_1 == 1'h0;
  assign _T_164 = _T_163 & valid_0;
  assign _T_165 = io_deq_ready ? valid_1 : _T_164;
  assign _T_166 = do_enq & _T_165;
  assign _T_167 = _T_160 | _T_166;
  assign _GEN_16 = _T_167 ? _T_156_btb_valid : elts_1_btb_valid;
  assign _GEN_18 = _T_167 ? _T_156_btb_bits_taken : elts_1_btb_bits_taken;
  assign _GEN_20 = _T_167 ? _T_156_btb_bits_bridx : elts_1_btb_bits_bridx;
  assign _GEN_26 = _T_167 ? _T_156_pc : elts_1_pc;
  assign _GEN_27 = _T_167 ? _T_156_data : elts_1_data;
  assign _GEN_29 = _T_167 ? _T_156_xcpt_pf_inst : elts_1_xcpt_pf_inst;
  assign _GEN_30 = _T_167 ? _T_156_xcpt_ae_inst : elts_1_xcpt_ae_inst;
  assign _GEN_31 = _T_167 ? _T_156_replay : elts_1_replay;
  assign _T_168_btb_valid = valid_3 ? elts_3_btb_valid : io_enq_bits_btb_valid;
  assign _T_168_btb_bits_taken = valid_3 ? elts_3_btb_bits_taken : io_enq_bits_btb_bits_taken;
  assign _T_168_btb_bits_bridx = valid_3 ? elts_3_btb_bits_bridx : io_enq_bits_btb_bits_bridx;
  assign _T_168_pc = valid_3 ? elts_3_pc : io_enq_bits_pc;
  assign _T_168_data = valid_3 ? elts_3_data : io_enq_bits_data;
  assign _T_168_xcpt_pf_inst = valid_3 ? elts_3_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst;
  assign _T_168_xcpt_ae_inst = valid_3 ? elts_3_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst;
  assign _T_168_replay = valid_3 ? elts_3_replay : io_enq_bits_replay;
  assign _T_172 = io_deq_ready & valid_3;
  assign _T_175 = valid_2 == 1'h0;
  assign _T_176 = _T_175 & valid_1;
  assign _T_177 = io_deq_ready ? valid_2 : _T_176;
  assign _T_178 = do_enq & _T_177;
  assign _T_179 = _T_172 | _T_178;
  assign _GEN_32 = _T_179 ? _T_168_btb_valid : elts_2_btb_valid;
  assign _GEN_34 = _T_179 ? _T_168_btb_bits_taken : elts_2_btb_bits_taken;
  assign _GEN_36 = _T_179 ? _T_168_btb_bits_bridx : elts_2_btb_bits_bridx;
  assign _GEN_42 = _T_179 ? _T_168_pc : elts_2_pc;
  assign _GEN_43 = _T_179 ? _T_168_data : elts_2_data;
  assign _GEN_45 = _T_179 ? _T_168_xcpt_pf_inst : elts_2_xcpt_pf_inst;
  assign _GEN_46 = _T_179 ? _T_168_xcpt_ae_inst : elts_2_xcpt_ae_inst;
  assign _GEN_47 = _T_179 ? _T_168_replay : elts_2_replay;
  assign _T_180_btb_valid = valid_4 ? elts_4_btb_valid : io_enq_bits_btb_valid;
  assign _T_180_btb_bits_taken = valid_4 ? elts_4_btb_bits_taken : io_enq_bits_btb_bits_taken;
  assign _T_180_btb_bits_bridx = valid_4 ? elts_4_btb_bits_bridx : io_enq_bits_btb_bits_bridx;
  assign _T_180_pc = valid_4 ? elts_4_pc : io_enq_bits_pc;
  assign _T_180_data = valid_4 ? elts_4_data : io_enq_bits_data;
  assign _T_180_xcpt_pf_inst = valid_4 ? elts_4_xcpt_pf_inst : io_enq_bits_xcpt_pf_inst;
  assign _T_180_xcpt_ae_inst = valid_4 ? elts_4_xcpt_ae_inst : io_enq_bits_xcpt_ae_inst;
  assign _T_180_replay = valid_4 ? elts_4_replay : io_enq_bits_replay;
  assign _T_184 = io_deq_ready & valid_4;
  assign _T_187 = valid_3 == 1'h0;
  assign _T_188 = _T_187 & valid_2;
  assign _T_189 = io_deq_ready ? valid_3 : _T_188;
  assign _T_190 = do_enq & _T_189;
  assign _T_191 = _T_184 | _T_190;
  assign _GEN_48 = _T_191 ? _T_180_btb_valid : elts_3_btb_valid;
  assign _GEN_50 = _T_191 ? _T_180_btb_bits_taken : elts_3_btb_bits_taken;
  assign _GEN_52 = _T_191 ? _T_180_btb_bits_bridx : elts_3_btb_bits_bridx;
  assign _GEN_58 = _T_191 ? _T_180_pc : elts_3_pc;
  assign _GEN_59 = _T_191 ? _T_180_data : elts_3_data;
  assign _GEN_61 = _T_191 ? _T_180_xcpt_pf_inst : elts_3_xcpt_pf_inst;
  assign _GEN_62 = _T_191 ? _T_180_xcpt_ae_inst : elts_3_xcpt_ae_inst;
  assign _GEN_63 = _T_191 ? _T_180_replay : elts_3_replay;
  assign _T_195 = valid_4 == 1'h0;
  assign _T_196 = _T_195 & valid_3;
  assign _T_197 = io_deq_ready ? valid_4 : _T_196;
  assign _T_198 = do_enq & _T_197;
  assign _GEN_64 = _T_198 ? io_enq_bits_btb_valid : elts_4_btb_valid;
  assign _GEN_66 = _T_198 ? io_enq_bits_btb_bits_taken : elts_4_btb_bits_taken;
  assign _GEN_68 = _T_198 ? io_enq_bits_btb_bits_bridx : elts_4_btb_bits_bridx;
  assign _GEN_74 = _T_198 ? io_enq_bits_pc : elts_4_pc;
  assign _GEN_75 = _T_198 ? io_enq_bits_data : elts_4_data;
  assign _GEN_77 = _T_198 ? io_enq_bits_xcpt_pf_inst : elts_4_xcpt_pf_inst;
  assign _GEN_78 = _T_198 ? io_enq_bits_xcpt_ae_inst : elts_4_xcpt_ae_inst;
  assign _GEN_79 = _T_198 ? io_enq_bits_replay : elts_4_replay;
  assign _T_201 = do_deq == 1'h0;
  assign _T_202 = do_enq & _T_201;
  assign _GEN_80 = _T_202 ? 1'h1 : valid_0;
  assign _T_206 = do_enq == 1'h0;
  assign _T_207 = _T_206 & do_deq;
  assign _T_210 = _T_207 & _T_163;
  assign _GEN_81 = _T_210 ? 1'h0 : _GEN_80;
  assign _T_215 = _T_202 & valid_0;
  assign _GEN_82 = _T_215 ? 1'h1 : valid_1;
  assign _T_222 = _T_207 & _T_175;
  assign _GEN_83 = _T_222 ? 1'h0 : _GEN_82;
  assign _T_227 = _T_202 & valid_1;
  assign _GEN_84 = _T_227 ? 1'h1 : valid_2;
  assign _T_234 = _T_207 & _T_187;
  assign _GEN_85 = _T_234 ? 1'h0 : _GEN_84;
  assign _T_239 = _T_202 & valid_2;
  assign _GEN_86 = _T_239 ? 1'h1 : valid_3;
  assign _T_246 = _T_207 & _T_195;
  assign _GEN_87 = _T_246 ? 1'h0 : _GEN_86;
  assign _T_251 = _T_202 & valid_3;
  assign _GEN_88 = _T_251 ? 1'h1 : valid_4;
  assign _GEN_89 = _T_207 ? 1'h0 : _GEN_88;
  assign _GEN_90 = io_enq_valid ? 1'h1 : valid_0;
  assign _GEN_91 = _T_150 ? io_enq_bits_btb_valid : elts_0_btb_valid;
  assign _GEN_93 = _T_150 ? io_enq_bits_btb_bits_taken : elts_0_btb_bits_taken;
  assign _GEN_95 = _T_150 ? io_enq_bits_btb_bits_bridx : elts_0_btb_bits_bridx;
  assign _GEN_101 = _T_150 ? io_enq_bits_pc : elts_0_pc;
  assign _GEN_102 = _T_150 ? io_enq_bits_data : elts_0_data;
  assign _GEN_104 = _T_150 ? io_enq_bits_xcpt_pf_inst : elts_0_xcpt_pf_inst;
  assign _GEN_105 = _T_150 ? io_enq_bits_xcpt_ae_inst : elts_0_xcpt_ae_inst;
  assign _GEN_106 = _T_150 ? io_enq_bits_replay : elts_0_replay;
  assign _T_265 = {valid_1,valid_0};
  assign _T_266 = {valid_4,valid_3};
  assign _T_267 = {_T_266,valid_2};
  assign _T_268 = {_T_267,_T_265};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  valid_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  valid_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  valid_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  valid_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  valid_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  elts_0_btb_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  elts_0_btb_bits_taken = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  elts_0_btb_bits_bridx = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  elts_0_pc = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  elts_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  elts_0_xcpt_pf_inst = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  elts_0_xcpt_ae_inst = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  elts_0_replay = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  elts_1_btb_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  elts_1_btb_bits_taken = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  elts_1_btb_bits_bridx = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  elts_1_pc = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  elts_1_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  elts_1_xcpt_pf_inst = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  elts_1_xcpt_ae_inst = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  elts_1_replay = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  elts_2_btb_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  elts_2_btb_bits_taken = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  elts_2_btb_bits_bridx = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  elts_2_pc = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  elts_2_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  elts_2_xcpt_pf_inst = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  elts_2_xcpt_ae_inst = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  elts_2_replay = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  elts_3_btb_valid = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  elts_3_btb_bits_taken = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  elts_3_btb_bits_bridx = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  elts_3_pc = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  elts_3_data = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  elts_3_xcpt_pf_inst = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  elts_3_xcpt_ae_inst = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  elts_3_replay = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  elts_4_btb_valid = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  elts_4_btb_bits_taken = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  elts_4_btb_bits_bridx = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  elts_4_pc = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  elts_4_data = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  elts_4_xcpt_pf_inst = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  elts_4_xcpt_ae_inst = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  elts_4_replay = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      valid_0 <= 1'h0;
    end else begin
      if (_T_210) begin
        valid_0 <= 1'h0;
      end else begin
        if (_T_202) begin
          valid_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      valid_1 <= 1'h0;
    end else begin
      if (_T_222) begin
        valid_1 <= 1'h0;
      end else begin
        if (_T_215) begin
          valid_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      valid_2 <= 1'h0;
    end else begin
      if (_T_234) begin
        valid_2 <= 1'h0;
      end else begin
        if (_T_227) begin
          valid_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      valid_3 <= 1'h0;
    end else begin
      if (_T_246) begin
        valid_3 <= 1'h0;
      end else begin
        if (_T_239) begin
          valid_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      valid_4 <= 1'h0;
    end else begin
      if (_T_207) begin
        valid_4 <= 1'h0;
      end else begin
        if (_T_251) begin
          valid_4 <= 1'h1;
        end
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_btb_valid <= elts_1_btb_valid;
      end else begin
        elts_0_btb_valid <= io_enq_bits_btb_valid;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_btb_bits_taken <= elts_1_btb_bits_taken;
      end else begin
        elts_0_btb_bits_taken <= io_enq_bits_btb_bits_taken;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_btb_bits_bridx <= elts_1_btb_bits_bridx;
      end else begin
        elts_0_btb_bits_bridx <= io_enq_bits_btb_bits_bridx;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_pc <= elts_1_pc;
      end else begin
        elts_0_pc <= io_enq_bits_pc;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_data <= elts_1_data;
      end else begin
        elts_0_data <= io_enq_bits_data;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_xcpt_pf_inst <= elts_1_xcpt_pf_inst;
      end else begin
        elts_0_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_xcpt_ae_inst <= elts_1_xcpt_ae_inst;
      end else begin
        elts_0_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (_T_155) begin
      if (valid_1) begin
        elts_0_replay <= elts_1_replay;
      end else begin
        elts_0_replay <= io_enq_bits_replay;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_btb_valid <= elts_2_btb_valid;
      end else begin
        elts_1_btb_valid <= io_enq_bits_btb_valid;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_btb_bits_taken <= elts_2_btb_bits_taken;
      end else begin
        elts_1_btb_bits_taken <= io_enq_bits_btb_bits_taken;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_btb_bits_bridx <= elts_2_btb_bits_bridx;
      end else begin
        elts_1_btb_bits_bridx <= io_enq_bits_btb_bits_bridx;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_pc <= elts_2_pc;
      end else begin
        elts_1_pc <= io_enq_bits_pc;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_data <= elts_2_data;
      end else begin
        elts_1_data <= io_enq_bits_data;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_xcpt_pf_inst <= elts_2_xcpt_pf_inst;
      end else begin
        elts_1_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_xcpt_ae_inst <= elts_2_xcpt_ae_inst;
      end else begin
        elts_1_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (_T_167) begin
      if (valid_2) begin
        elts_1_replay <= elts_2_replay;
      end else begin
        elts_1_replay <= io_enq_bits_replay;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_btb_valid <= elts_3_btb_valid;
      end else begin
        elts_2_btb_valid <= io_enq_bits_btb_valid;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_btb_bits_taken <= elts_3_btb_bits_taken;
      end else begin
        elts_2_btb_bits_taken <= io_enq_bits_btb_bits_taken;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_btb_bits_bridx <= elts_3_btb_bits_bridx;
      end else begin
        elts_2_btb_bits_bridx <= io_enq_bits_btb_bits_bridx;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_pc <= elts_3_pc;
      end else begin
        elts_2_pc <= io_enq_bits_pc;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_data <= elts_3_data;
      end else begin
        elts_2_data <= io_enq_bits_data;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_xcpt_pf_inst <= elts_3_xcpt_pf_inst;
      end else begin
        elts_2_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_xcpt_ae_inst <= elts_3_xcpt_ae_inst;
      end else begin
        elts_2_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (_T_179) begin
      if (valid_3) begin
        elts_2_replay <= elts_3_replay;
      end else begin
        elts_2_replay <= io_enq_bits_replay;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_btb_valid <= elts_4_btb_valid;
      end else begin
        elts_3_btb_valid <= io_enq_bits_btb_valid;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_btb_bits_taken <= elts_4_btb_bits_taken;
      end else begin
        elts_3_btb_bits_taken <= io_enq_bits_btb_bits_taken;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_btb_bits_bridx <= elts_4_btb_bits_bridx;
      end else begin
        elts_3_btb_bits_bridx <= io_enq_bits_btb_bits_bridx;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_pc <= elts_4_pc;
      end else begin
        elts_3_pc <= io_enq_bits_pc;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_data <= elts_4_data;
      end else begin
        elts_3_data <= io_enq_bits_data;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_xcpt_pf_inst <= elts_4_xcpt_pf_inst;
      end else begin
        elts_3_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_xcpt_ae_inst <= elts_4_xcpt_ae_inst;
      end else begin
        elts_3_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
      end
    end
    if (_T_191) begin
      if (valid_4) begin
        elts_3_replay <= elts_4_replay;
      end else begin
        elts_3_replay <= io_enq_bits_replay;
      end
    end
    if (_T_198) begin
      elts_4_btb_valid <= io_enq_bits_btb_valid;
    end
    if (_T_198) begin
      elts_4_btb_bits_taken <= io_enq_bits_btb_bits_taken;
    end
    if (_T_198) begin
      elts_4_btb_bits_bridx <= io_enq_bits_btb_bits_bridx;
    end
    if (_T_198) begin
      elts_4_pc <= io_enq_bits_pc;
    end
    if (_T_198) begin
      elts_4_data <= io_enq_bits_data;
    end
    if (_T_198) begin
      elts_4_xcpt_pf_inst <= io_enq_bits_xcpt_pf_inst;
    end
    if (_T_198) begin
      elts_4_xcpt_ae_inst <= io_enq_bits_xcpt_ae_inst;
    end
    if (_T_198) begin
      elts_4_replay <= io_enq_bits_replay;
    end
  end
endmodule
module Frontend_frontend(
  input         clock,
  input         reset,
  input         io_tl_out_0_a_ready,
  output        io_tl_out_0_a_valid,
  output [2:0]  io_tl_out_0_a_bits_opcode,
  output [2:0]  io_tl_out_0_a_bits_param,
  output [3:0]  io_tl_out_0_a_bits_size,
  output        io_tl_out_0_a_bits_source,
  output [31:0] io_tl_out_0_a_bits_address,
  output [3:0]  io_tl_out_0_a_bits_mask,
  output [31:0] io_tl_out_0_a_bits_data,
  output        io_tl_out_0_d_ready,
  input         io_tl_out_0_d_valid,
  input  [2:0]  io_tl_out_0_d_bits_opcode,
  input  [3:0]  io_tl_out_0_d_bits_size,
  input  [31:0] io_tl_out_0_d_bits_data,
  input         io_tl_out_0_d_bits_error,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_pc,
  input         io_cpu_req_bits_speculative,
  input         io_cpu_resp_ready,
  output        io_cpu_resp_valid,
  output        io_cpu_resp_bits_btb_valid,
  output        io_cpu_resp_bits_btb_bits_taken,
  output        io_cpu_resp_bits_btb_bits_bridx,
  output [31:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cpu_resp_bits_xcpt_pf_inst,
  output        io_cpu_resp_bits_xcpt_ae_inst,
  output        io_cpu_resp_bits_replay,
  input         io_cpu_flush_icache,
  output [31:0] io_cpu_npc,
  output        io_ptw_req_valid,
  output [19:0] io_ptw_req_bits_addr,
  input         io_ptw_resp_valid,
  input  [1:0]  io_ptw_status_dprv,
  input  [1:0]  io_ptw_status_prv,
  input         io_ptw_status_mxr,
  input         io_ptw_status_sum,
  input         io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
  input         io_ptw_pmp_0_cfg_w,
  input         io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
  input         io_ptw_pmp_1_cfg_w,
  input         io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
  input         io_ptw_pmp_2_cfg_w,
  input         io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
  input         io_ptw_pmp_3_cfg_w,
  input         io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
  input         io_ptw_pmp_4_cfg_w,
  input         io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
  input         io_ptw_pmp_5_cfg_w,
  input         io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
  input         io_ptw_pmp_6_cfg_w,
  input         io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
  input         io_ptw_pmp_7_cfg_w,
  input         io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input  [31:0] io_resetVector
);
  wire  icache_clock;
  wire  icache_reset;
  wire  icache_io_req_ready;
  wire  icache_io_req_valid;
  wire [31:0] icache_io_req_bits_addr;
  wire [31:0] icache_io_s1_paddr;
  wire  icache_io_s1_kill;
  wire  icache_io_s2_kill;
  wire  icache_io_resp_valid;
  wire [31:0] icache_io_resp_bits_data;
  wire  icache_io_resp_bits_ae;
  wire  icache_io_invalidate;
  wire  icache_io_tl_out_0_a_ready;
  wire  icache_io_tl_out_0_a_valid;
  wire [2:0] icache_io_tl_out_0_a_bits_opcode;
  wire [2:0] icache_io_tl_out_0_a_bits_param;
  wire [3:0] icache_io_tl_out_0_a_bits_size;
  wire  icache_io_tl_out_0_a_bits_source;
  wire [31:0] icache_io_tl_out_0_a_bits_address;
  wire [3:0] icache_io_tl_out_0_a_bits_mask;
  wire [31:0] icache_io_tl_out_0_a_bits_data;
  wire  icache_io_tl_out_0_d_ready;
  wire  icache_io_tl_out_0_d_valid;
  wire [2:0] icache_io_tl_out_0_d_bits_opcode;
  wire [3:0] icache_io_tl_out_0_d_bits_size;
  wire [31:0] icache_io_tl_out_0_d_bits_data;
  wire  icache_io_tl_out_0_d_bits_error;
  wire  tlb_clock;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [31:0] tlb_io_req_bits_vaddr;
  wire  tlb_io_req_bits_instruction;
  wire [1:0] tlb_io_req_bits_size;
  wire [4:0] tlb_io_req_bits_cmd;
  wire  tlb_io_resp_miss;
  wire [31:0] tlb_io_resp_paddr;
  wire  tlb_io_resp_pf_ld;
  wire  tlb_io_resp_pf_st;
  wire  tlb_io_resp_pf_inst;
  wire  tlb_io_resp_ae_ld;
  wire  tlb_io_resp_ae_st;
  wire  tlb_io_resp_ae_inst;
  wire  tlb_io_resp_ma_ld;
  wire  tlb_io_resp_ma_st;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_valid;
  wire [19:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_resp_valid;
  wire [1:0] tlb_io_ptw_status_dprv;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_sum;
  wire  tlb_io_ptw_pmp_0_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_0_cfg_a;
  wire  tlb_io_ptw_pmp_0_cfg_x;
  wire  tlb_io_ptw_pmp_0_cfg_w;
  wire  tlb_io_ptw_pmp_0_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_0_addr;
  wire [31:0] tlb_io_ptw_pmp_0_mask;
  wire  tlb_io_ptw_pmp_1_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_1_cfg_a;
  wire  tlb_io_ptw_pmp_1_cfg_x;
  wire  tlb_io_ptw_pmp_1_cfg_w;
  wire  tlb_io_ptw_pmp_1_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_1_addr;
  wire [31:0] tlb_io_ptw_pmp_1_mask;
  wire  tlb_io_ptw_pmp_2_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_2_cfg_a;
  wire  tlb_io_ptw_pmp_2_cfg_x;
  wire  tlb_io_ptw_pmp_2_cfg_w;
  wire  tlb_io_ptw_pmp_2_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_2_addr;
  wire [31:0] tlb_io_ptw_pmp_2_mask;
  wire  tlb_io_ptw_pmp_3_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_3_cfg_a;
  wire  tlb_io_ptw_pmp_3_cfg_x;
  wire  tlb_io_ptw_pmp_3_cfg_w;
  wire  tlb_io_ptw_pmp_3_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_3_addr;
  wire [31:0] tlb_io_ptw_pmp_3_mask;
  wire  tlb_io_ptw_pmp_4_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_4_cfg_a;
  wire  tlb_io_ptw_pmp_4_cfg_x;
  wire  tlb_io_ptw_pmp_4_cfg_w;
  wire  tlb_io_ptw_pmp_4_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_4_addr;
  wire [31:0] tlb_io_ptw_pmp_4_mask;
  wire  tlb_io_ptw_pmp_5_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_5_cfg_a;
  wire  tlb_io_ptw_pmp_5_cfg_x;
  wire  tlb_io_ptw_pmp_5_cfg_w;
  wire  tlb_io_ptw_pmp_5_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_5_addr;
  wire [31:0] tlb_io_ptw_pmp_5_mask;
  wire  tlb_io_ptw_pmp_6_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_6_cfg_a;
  wire  tlb_io_ptw_pmp_6_cfg_x;
  wire  tlb_io_ptw_pmp_6_cfg_w;
  wire  tlb_io_ptw_pmp_6_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_6_addr;
  wire [31:0] tlb_io_ptw_pmp_6_mask;
  wire  tlb_io_ptw_pmp_7_cfg_l;
  wire [1:0] tlb_io_ptw_pmp_7_cfg_a;
  wire  tlb_io_ptw_pmp_7_cfg_x;
  wire  tlb_io_ptw_pmp_7_cfg_w;
  wire  tlb_io_ptw_pmp_7_cfg_r;
  wire [29:0] tlb_io_ptw_pmp_7_addr;
  wire [31:0] tlb_io_ptw_pmp_7_mask;
  wire  _T_197;
  wire  fq_clock;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire  fq_io_enq_bits_btb_valid;
  wire  fq_io_enq_bits_btb_bits_taken;
  wire  fq_io_enq_bits_btb_bits_bridx;
  wire [31:0] fq_io_enq_bits_pc;
  wire [31:0] fq_io_enq_bits_data;
  wire  fq_io_enq_bits_xcpt_pf_inst;
  wire  fq_io_enq_bits_xcpt_ae_inst;
  wire  fq_io_enq_bits_replay;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire  fq_io_deq_bits_btb_valid;
  wire  fq_io_deq_bits_btb_bits_taken;
  wire  fq_io_deq_bits_btb_bits_bridx;
  wire [31:0] fq_io_deq_bits_pc;
  wire [31:0] fq_io_deq_bits_data;
  wire  fq_io_deq_bits_xcpt_pf_inst;
  wire  fq_io_deq_bits_xcpt_ae_inst;
  wire  fq_io_deq_bits_replay;
  wire [4:0] fq_io_mask;
  wire  _T_202;
  wire  _T_204;
  wire  s0_valid;
  reg [31:0] s1_pc;
  reg [31:0] _RAND_0;
  reg  s1_speculative;
  reg [31:0] _RAND_1;
  reg  s2_valid;
  reg [31:0] _RAND_2;
  wire [31:0] _T_209;
  wire [31:0] _T_211;
  wire [31:0] _T_212;
  reg [31:0] s2_pc;
  reg [31:0] _RAND_3;
  reg  s2_btb_resp_bits_taken;
  reg [31:0] _RAND_4;
  reg  s2_btb_resp_bits_bridx;
  reg [31:0] _RAND_5;
  reg  s2_tlb_resp_miss;
  reg [31:0] _RAND_6;
  reg  s2_tlb_resp_pf_inst;
  reg [31:0] _RAND_7;
  reg  s2_tlb_resp_ae_inst;
  reg [31:0] _RAND_8;
  reg  s2_tlb_resp_cacheable;
  reg [31:0] _RAND_9;
  wire  _T_216;
  wire [1:0] _T_217;
  wire  _T_219;
  wire  s2_xcpt;
  reg  s2_speculative;
  reg [31:0] _RAND_10;
  wire [31:0] _T_226;
  wire [31:0] _T_228;
  wire [31:0] s1_base_pc;
  wire [32:0] _T_230;
  wire [31:0] ntpc;
  wire  _T_235;
  wire  _T_237;
  wire  _T_238;
  wire  _T_240;
  wire  _T_241;
  reg  _T_244;
  reg [31:0] _RAND_11;
  wire  _T_245;
  wire [31:0] npc;
  wire  _T_247;
  wire  _T_248;
  wire  _T_249;
  wire  _T_250;
  wire  _T_251;
  wire  _T_255;
  wire  _T_257;
  wire  _T_258;
  wire [31:0] _GEN_1;
  wire  _GEN_2;
  wire  _GEN_3;
  wire  _GEN_7;
  wire  _GEN_10;
  wire  _GEN_14;
  wire  _T_265;
  wire  _T_266;
  wire  _T_268;
  wire  _T_269;
  wire  _T_270;
  wire  _T_271;
  wire  _T_272;
  wire  _T_273;
  wire [31:0] _T_274;
  wire [31:0] _T_275;
  wire [31:0] _T_277;
  wire [31:0] _T_278;
  wire  _T_283;
  wire  _T_284;
  wire  _T_286;
  wire  _T_287;
  wire  _T_288;
  wire  _GEN_15;
  ICache_icache icache (
    .clock(icache_clock),
    .reset(icache_reset),
    .io_req_ready(icache_io_req_ready),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_paddr(icache_io_s1_paddr),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_ae(icache_io_resp_bits_ae),
    .io_invalidate(icache_io_invalidate),
    .io_tl_out_0_a_ready(icache_io_tl_out_0_a_ready),
    .io_tl_out_0_a_valid(icache_io_tl_out_0_a_valid),
    .io_tl_out_0_a_bits_opcode(icache_io_tl_out_0_a_bits_opcode),
    .io_tl_out_0_a_bits_param(icache_io_tl_out_0_a_bits_param),
    .io_tl_out_0_a_bits_size(icache_io_tl_out_0_a_bits_size),
    .io_tl_out_0_a_bits_source(icache_io_tl_out_0_a_bits_source),
    .io_tl_out_0_a_bits_address(icache_io_tl_out_0_a_bits_address),
    .io_tl_out_0_a_bits_mask(icache_io_tl_out_0_a_bits_mask),
    .io_tl_out_0_a_bits_data(icache_io_tl_out_0_a_bits_data),
    .io_tl_out_0_d_ready(icache_io_tl_out_0_d_ready),
    .io_tl_out_0_d_valid(icache_io_tl_out_0_d_valid),
    .io_tl_out_0_d_bits_opcode(icache_io_tl_out_0_d_bits_opcode),
    .io_tl_out_0_d_bits_size(icache_io_tl_out_0_d_bits_size),
    .io_tl_out_0_d_bits_data(icache_io_tl_out_0_d_bits_data),
    .io_tl_out_0_d_bits_error(icache_io_tl_out_0_d_bits_error)
  );
  TLB tlb (
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vaddr(tlb_io_req_bits_vaddr),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_size(tlb_io_req_bits_size),
    .io_req_bits_cmd(tlb_io_req_bits_cmd),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_paddr(tlb_io_resp_paddr),
    .io_resp_pf_ld(tlb_io_resp_pf_ld),
    .io_resp_pf_st(tlb_io_resp_pf_st),
    .io_resp_pf_inst(tlb_io_resp_pf_inst),
    .io_resp_ae_ld(tlb_io_resp_ae_ld),
    .io_resp_ae_st(tlb_io_resp_ae_st),
    .io_resp_ae_inst(tlb_io_resp_ae_inst),
    .io_resp_ma_ld(tlb_io_resp_ma_ld),
    .io_resp_ma_st(tlb_io_resp_ma_st),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_status_dprv(tlb_io_ptw_status_dprv),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_sum(tlb_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(tlb_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(tlb_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(tlb_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(tlb_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(tlb_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(tlb_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(tlb_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(tlb_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(tlb_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(tlb_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(tlb_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(tlb_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(tlb_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(tlb_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(tlb_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(tlb_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(tlb_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(tlb_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(tlb_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(tlb_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(tlb_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(tlb_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(tlb_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(tlb_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(tlb_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(tlb_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(tlb_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(tlb_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(tlb_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(tlb_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(tlb_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(tlb_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(tlb_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(tlb_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(tlb_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(tlb_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(tlb_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(tlb_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(tlb_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(tlb_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(tlb_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(tlb_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(tlb_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(tlb_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(tlb_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(tlb_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(tlb_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(tlb_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(tlb_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(tlb_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(tlb_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(tlb_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(tlb_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(tlb_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(tlb_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(tlb_io_ptw_pmp_7_mask)
  );
  ShiftQueue fq (
    .clock(fq_clock),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_btb_valid(fq_io_enq_bits_btb_valid),
    .io_enq_bits_btb_bits_taken(fq_io_enq_bits_btb_bits_taken),
    .io_enq_bits_btb_bits_bridx(fq_io_enq_bits_btb_bits_bridx),
    .io_enq_bits_pc(fq_io_enq_bits_pc),
    .io_enq_bits_data(fq_io_enq_bits_data),
    .io_enq_bits_xcpt_pf_inst(fq_io_enq_bits_xcpt_pf_inst),
    .io_enq_bits_xcpt_ae_inst(fq_io_enq_bits_xcpt_ae_inst),
    .io_enq_bits_replay(fq_io_enq_bits_replay),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_btb_valid(fq_io_deq_bits_btb_valid),
    .io_deq_bits_btb_bits_taken(fq_io_deq_bits_btb_bits_taken),
    .io_deq_bits_btb_bits_bridx(fq_io_deq_bits_btb_bits_bridx),
    .io_deq_bits_pc(fq_io_deq_bits_pc),
    .io_deq_bits_data(fq_io_deq_bits_data),
    .io_deq_bits_xcpt_pf_inst(fq_io_deq_bits_xcpt_pf_inst),
    .io_deq_bits_xcpt_ae_inst(fq_io_deq_bits_xcpt_ae_inst),
    .io_deq_bits_replay(fq_io_deq_bits_replay),
    .io_mask(fq_io_mask)
  );
  assign io_tl_out_0_a_valid = icache_io_tl_out_0_a_valid;
  assign io_tl_out_0_a_bits_opcode = icache_io_tl_out_0_a_bits_opcode;
  assign io_tl_out_0_a_bits_param = icache_io_tl_out_0_a_bits_param;
  assign io_tl_out_0_a_bits_size = icache_io_tl_out_0_a_bits_size;
  assign io_tl_out_0_a_bits_source = icache_io_tl_out_0_a_bits_source;
  assign io_tl_out_0_a_bits_address = icache_io_tl_out_0_a_bits_address;
  assign io_tl_out_0_a_bits_mask = icache_io_tl_out_0_a_bits_mask;
  assign io_tl_out_0_a_bits_data = icache_io_tl_out_0_a_bits_data;
  assign io_tl_out_0_d_ready = icache_io_tl_out_0_d_ready;
  assign io_cpu_resp_valid = fq_io_deq_valid;
  assign io_cpu_resp_bits_btb_valid = fq_io_deq_bits_btb_valid;
  assign io_cpu_resp_bits_btb_bits_taken = fq_io_deq_bits_btb_bits_taken;
  assign io_cpu_resp_bits_btb_bits_bridx = fq_io_deq_bits_btb_bits_bridx;
  assign io_cpu_resp_bits_pc = fq_io_deq_bits_pc;
  assign io_cpu_resp_bits_data = fq_io_deq_bits_data;
  assign io_cpu_resp_bits_xcpt_pf_inst = fq_io_deq_bits_xcpt_pf_inst;
  assign io_cpu_resp_bits_xcpt_ae_inst = fq_io_deq_bits_xcpt_ae_inst;
  assign io_cpu_resp_bits_replay = fq_io_deq_bits_replay;
  assign io_cpu_npc = _T_278;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_req_valid = s0_valid;
  assign icache_io_req_bits_addr = io_cpu_npc;
  assign icache_io_s1_paddr = tlb_io_resp_paddr;
  assign icache_io_s1_kill = _T_266;
  assign icache_io_s2_kill = _T_271;
  assign icache_io_invalidate = io_cpu_flush_icache;
  assign icache_io_tl_out_0_a_ready = io_tl_out_0_a_ready;
  assign icache_io_tl_out_0_d_valid = io_tl_out_0_d_valid;
  assign icache_io_tl_out_0_d_bits_opcode = io_tl_out_0_d_bits_opcode;
  assign icache_io_tl_out_0_d_bits_size = io_tl_out_0_d_bits_size;
  assign icache_io_tl_out_0_d_bits_data = io_tl_out_0_d_bits_data;
  assign icache_io_tl_out_0_d_bits_error = io_tl_out_0_d_bits_error;
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = _T_255;
  assign tlb_io_req_bits_vaddr = s1_pc;
  assign tlb_io_req_bits_instruction = 1'h1;
  assign tlb_io_req_bits_size = 2'h2;
  assign tlb_io_req_bits_cmd = 5'h0;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_status_dprv = io_ptw_status_dprv;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_sum = io_ptw_status_sum;
  assign tlb_io_ptw_pmp_0_cfg_l = io_ptw_pmp_0_cfg_l;
  assign tlb_io_ptw_pmp_0_cfg_a = io_ptw_pmp_0_cfg_a;
  assign tlb_io_ptw_pmp_0_cfg_x = io_ptw_pmp_0_cfg_x;
  assign tlb_io_ptw_pmp_0_cfg_w = io_ptw_pmp_0_cfg_w;
  assign tlb_io_ptw_pmp_0_cfg_r = io_ptw_pmp_0_cfg_r;
  assign tlb_io_ptw_pmp_0_addr = io_ptw_pmp_0_addr;
  assign tlb_io_ptw_pmp_0_mask = io_ptw_pmp_0_mask;
  assign tlb_io_ptw_pmp_1_cfg_l = io_ptw_pmp_1_cfg_l;
  assign tlb_io_ptw_pmp_1_cfg_a = io_ptw_pmp_1_cfg_a;
  assign tlb_io_ptw_pmp_1_cfg_x = io_ptw_pmp_1_cfg_x;
  assign tlb_io_ptw_pmp_1_cfg_w = io_ptw_pmp_1_cfg_w;
  assign tlb_io_ptw_pmp_1_cfg_r = io_ptw_pmp_1_cfg_r;
  assign tlb_io_ptw_pmp_1_addr = io_ptw_pmp_1_addr;
  assign tlb_io_ptw_pmp_1_mask = io_ptw_pmp_1_mask;
  assign tlb_io_ptw_pmp_2_cfg_l = io_ptw_pmp_2_cfg_l;
  assign tlb_io_ptw_pmp_2_cfg_a = io_ptw_pmp_2_cfg_a;
  assign tlb_io_ptw_pmp_2_cfg_x = io_ptw_pmp_2_cfg_x;
  assign tlb_io_ptw_pmp_2_cfg_w = io_ptw_pmp_2_cfg_w;
  assign tlb_io_ptw_pmp_2_cfg_r = io_ptw_pmp_2_cfg_r;
  assign tlb_io_ptw_pmp_2_addr = io_ptw_pmp_2_addr;
  assign tlb_io_ptw_pmp_2_mask = io_ptw_pmp_2_mask;
  assign tlb_io_ptw_pmp_3_cfg_l = io_ptw_pmp_3_cfg_l;
  assign tlb_io_ptw_pmp_3_cfg_a = io_ptw_pmp_3_cfg_a;
  assign tlb_io_ptw_pmp_3_cfg_x = io_ptw_pmp_3_cfg_x;
  assign tlb_io_ptw_pmp_3_cfg_w = io_ptw_pmp_3_cfg_w;
  assign tlb_io_ptw_pmp_3_cfg_r = io_ptw_pmp_3_cfg_r;
  assign tlb_io_ptw_pmp_3_addr = io_ptw_pmp_3_addr;
  assign tlb_io_ptw_pmp_3_mask = io_ptw_pmp_3_mask;
  assign tlb_io_ptw_pmp_4_cfg_l = io_ptw_pmp_4_cfg_l;
  assign tlb_io_ptw_pmp_4_cfg_a = io_ptw_pmp_4_cfg_a;
  assign tlb_io_ptw_pmp_4_cfg_x = io_ptw_pmp_4_cfg_x;
  assign tlb_io_ptw_pmp_4_cfg_w = io_ptw_pmp_4_cfg_w;
  assign tlb_io_ptw_pmp_4_cfg_r = io_ptw_pmp_4_cfg_r;
  assign tlb_io_ptw_pmp_4_addr = io_ptw_pmp_4_addr;
  assign tlb_io_ptw_pmp_4_mask = io_ptw_pmp_4_mask;
  assign tlb_io_ptw_pmp_5_cfg_l = io_ptw_pmp_5_cfg_l;
  assign tlb_io_ptw_pmp_5_cfg_a = io_ptw_pmp_5_cfg_a;
  assign tlb_io_ptw_pmp_5_cfg_x = io_ptw_pmp_5_cfg_x;
  assign tlb_io_ptw_pmp_5_cfg_w = io_ptw_pmp_5_cfg_w;
  assign tlb_io_ptw_pmp_5_cfg_r = io_ptw_pmp_5_cfg_r;
  assign tlb_io_ptw_pmp_5_addr = io_ptw_pmp_5_addr;
  assign tlb_io_ptw_pmp_5_mask = io_ptw_pmp_5_mask;
  assign tlb_io_ptw_pmp_6_cfg_l = io_ptw_pmp_6_cfg_l;
  assign tlb_io_ptw_pmp_6_cfg_a = io_ptw_pmp_6_cfg_a;
  assign tlb_io_ptw_pmp_6_cfg_x = io_ptw_pmp_6_cfg_x;
  assign tlb_io_ptw_pmp_6_cfg_w = io_ptw_pmp_6_cfg_w;
  assign tlb_io_ptw_pmp_6_cfg_r = io_ptw_pmp_6_cfg_r;
  assign tlb_io_ptw_pmp_6_addr = io_ptw_pmp_6_addr;
  assign tlb_io_ptw_pmp_6_mask = io_ptw_pmp_6_mask;
  assign tlb_io_ptw_pmp_7_cfg_l = io_ptw_pmp_7_cfg_l;
  assign tlb_io_ptw_pmp_7_cfg_a = io_ptw_pmp_7_cfg_a;
  assign tlb_io_ptw_pmp_7_cfg_x = io_ptw_pmp_7_cfg_x;
  assign tlb_io_ptw_pmp_7_cfg_w = io_ptw_pmp_7_cfg_w;
  assign tlb_io_ptw_pmp_7_cfg_r = io_ptw_pmp_7_cfg_r;
  assign tlb_io_ptw_pmp_7_addr = io_ptw_pmp_7_addr;
  assign tlb_io_ptw_pmp_7_mask = io_ptw_pmp_7_mask;
  assign _T_197 = reset | io_cpu_req_valid;
  assign fq_clock = clock;
  assign fq_reset = _T_197;
  assign fq_io_enq_valid = _T_273;
  assign fq_io_enq_bits_btb_valid = 1'h0;
  assign fq_io_enq_bits_btb_bits_taken = s2_btb_resp_bits_taken;
  assign fq_io_enq_bits_btb_bits_bridx = s2_btb_resp_bits_bridx;
  assign fq_io_enq_bits_pc = s2_pc;
  assign fq_io_enq_bits_data = icache_io_resp_bits_data;
  assign fq_io_enq_bits_xcpt_pf_inst = s2_tlb_resp_pf_inst;
  assign fq_io_enq_bits_xcpt_ae_inst = _GEN_15;
  assign fq_io_enq_bits_replay = _T_287;
  assign fq_io_deq_ready = io_cpu_resp_ready;
  assign _T_202 = fq_io_mask[2];
  assign _T_204 = _T_202 == 1'h0;
  assign s0_valid = io_cpu_req_valid | _T_204;
  assign _T_209 = ~ io_resetVector;
  assign _T_211 = _T_209 | 32'h1;
  assign _T_212 = ~ _T_211;
  assign _T_216 = s2_tlb_resp_miss == 1'h0;
  assign _T_217 = {fq_io_enq_bits_xcpt_pf_inst,fq_io_enq_bits_xcpt_ae_inst};
  assign _T_219 = _T_217 != 2'h0;
  assign s2_xcpt = _T_216 & _T_219;
  assign _T_226 = ~ s1_pc;
  assign _T_228 = _T_226 | 32'h3;
  assign s1_base_pc = ~ _T_228;
  assign _T_230 = s1_base_pc + 32'h4;
  assign ntpc = _T_230[31:0];
  assign _T_235 = fq_io_enq_ready & fq_io_enq_valid;
  assign _T_237 = _T_235 == 1'h0;
  assign _T_238 = s2_valid & _T_237;
  assign _T_240 = s0_valid == 1'h0;
  assign _T_241 = _T_245 & _T_240;
  assign _T_245 = _T_238 | _T_244;
  assign npc = _T_245 ? s2_pc : ntpc;
  assign _T_247 = s2_speculative == 1'h0;
  assign _T_248 = s2_valid & _T_247;
  assign _T_249 = s1_speculative | _T_248;
  assign _T_250 = _T_245 ? s2_speculative : _T_249;
  assign _T_251 = io_cpu_req_valid ? io_cpu_req_bits_speculative : _T_250;
  assign _T_255 = _T_245 == 1'h0;
  assign _T_257 = io_cpu_req_valid == 1'h0;
  assign _T_258 = _T_255 & _T_257;
  assign _GEN_1 = _T_258 ? s1_pc : s2_pc;
  assign _GEN_2 = _T_258 ? s1_speculative : s2_speculative;
  assign _GEN_3 = _T_258 ? tlb_io_resp_miss : s2_tlb_resp_miss;
  assign _GEN_7 = _T_258 ? tlb_io_resp_pf_inst : s2_tlb_resp_pf_inst;
  assign _GEN_10 = _T_258 ? tlb_io_resp_ae_inst : s2_tlb_resp_ae_inst;
  assign _GEN_14 = _T_258 ? tlb_io_resp_cacheable : s2_tlb_resp_cacheable;
  assign _T_265 = io_cpu_req_valid | tlb_io_resp_miss;
  assign _T_266 = _T_265 | _T_245;
  assign _T_268 = s2_tlb_resp_cacheable == 1'h0;
  assign _T_269 = s2_speculative & _T_268;
  assign _T_270 = _T_269 | s2_xcpt;
  assign _T_271 = s2_valid & _T_270;
  assign _T_272 = icache_io_resp_valid | icache_io_s2_kill;
  assign _T_273 = s2_valid & _T_272;
  assign _T_274 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign _T_275 = ~ _T_274;
  assign _T_277 = _T_275 | 32'h1;
  assign _T_278 = ~ _T_277;
  assign _T_283 = icache_io_resp_valid == 1'h0;
  assign _T_284 = icache_io_s2_kill & _T_283;
  assign _T_286 = s2_xcpt == 1'h0;
  assign _T_287 = _T_284 & _T_286;
  assign _T_288 = icache_io_resp_valid & icache_io_resp_bits_ae;
  assign _GEN_15 = _T_288 ? 1'h1 : s2_tlb_resp_ae_inst;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  s1_pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  s1_speculative = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  s2_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  s2_pc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  s2_btb_resp_bits_taken = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  s2_btb_resp_bits_bridx = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  s2_tlb_resp_miss = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  s2_tlb_resp_pf_inst = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  s2_tlb_resp_ae_inst = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  s2_tlb_resp_cacheable = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  s2_speculative = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_244 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    s1_pc <= io_cpu_npc;
    if (io_cpu_req_valid) begin
      s1_speculative <= io_cpu_req_bits_speculative;
    end else begin
      if (_T_245) begin
        s1_speculative <= s2_speculative;
      end else begin
        s1_speculative <= _T_249;
      end
    end
    if (reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= _T_258;
    end
    if (reset) begin
      s2_pc <= _T_212;
    end else begin
      if (_T_258) begin
        s2_pc <= s1_pc;
      end
    end
    if (_T_258) begin
      s2_tlb_resp_miss <= tlb_io_resp_miss;
    end
    if (_T_258) begin
      s2_tlb_resp_pf_inst <= tlb_io_resp_pf_inst;
    end
    if (_T_258) begin
      s2_tlb_resp_ae_inst <= tlb_io_resp_ae_inst;
    end
    if (_T_258) begin
      s2_tlb_resp_cacheable <= tlb_io_resp_cacheable;
    end
    if (reset) begin
      s2_speculative <= 1'h0;
    end else begin
      if (_T_258) begin
        s2_speculative <= s1_speculative;
      end
    end
    if (reset) begin
      _T_244 <= 1'h1;
    end else begin
      _T_244 <= _T_241;
    end
  end
endmodule
module ScratchpadSlavePort(
  input         clock,
  input         reset,
  output        io_tl_in_0_a_ready,
  input         io_tl_in_0_a_valid,
  input  [2:0]  io_tl_in_0_a_bits_opcode,
  input  [2:0]  io_tl_in_0_a_bits_param,
  input  [1:0]  io_tl_in_0_a_bits_size,
  input  [9:0]  io_tl_in_0_a_bits_source,
  input  [31:0] io_tl_in_0_a_bits_address,
  input  [3:0]  io_tl_in_0_a_bits_mask,
  input  [31:0] io_tl_in_0_a_bits_data,
  input         io_tl_in_0_d_ready,
  output        io_tl_in_0_d_valid,
  output [2:0]  io_tl_in_0_d_bits_opcode,
  output [1:0]  io_tl_in_0_d_bits_param,
  output [1:0]  io_tl_in_0_d_bits_size,
  output [9:0]  io_tl_in_0_d_bits_source,
  output        io_tl_in_0_d_bits_sink,
  output [31:0] io_tl_in_0_d_bits_data,
  output        io_tl_in_0_d_bits_error,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [2:0]  io_dmem_req_bits_typ,
  output        io_dmem_req_bits_phys,
  output        io_dmem_s1_kill,
  output [31:0] io_dmem_s1_data_data,
  output [3:0]  io_dmem_s1_data_mask,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [31:0] io_dmem_resp_bits_data_raw,
  output        io_dmem_invalidate_lr
);
  reg [1:0] state;
  reg [31:0] _RAND_0;
  wire [1:0] _GEN_0;
  wire  _T_80;
  wire [1:0] _GEN_1;
  wire [1:0] _GEN_2;
  wire  _T_81;
  wire [1:0] _GEN_3;
  reg [2:0] acq_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] acq_param;
  reg [31:0] _RAND_2;
  reg [1:0] acq_size;
  reg [31:0] _RAND_3;
  reg [9:0] acq_source;
  reg [31:0] _RAND_4;
  reg [31:0] acq_address;
  reg [31:0] _RAND_5;
  reg [3:0] acq_mask;
  reg [31:0] _RAND_6;
  reg [31:0] acq_data;
  reg [31:0] _RAND_7;
  wire [31:0] _GEN_4;
  wire  _T_82;
  wire [2:0] _GEN_5;
  wire [2:0] _GEN_6;
  wire [1:0] _GEN_7;
  wire [9:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [3:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire  _T_83;
  wire  ready;
  wire  _T_85;
  wire  _T_86;
  wire  _T_87;
  wire  _T_88;
  wire [2:0] _T_90_opcode;
  wire [2:0] _T_90_param;
  wire [1:0] _T_90_size;
  wire [31:0] _T_90_address;
  wire [2:0] _T_92_typ;
  wire  _T_112;
  wire [3:0] _T_113;
  wire  _T_114;
  wire [3:0] _T_115;
  wire  _T_116;
  wire [3:0] _T_117;
  wire  _T_118;
  wire [3:0] _T_119;
  wire  _T_120;
  wire [3:0] _T_121;
  wire [2:0] _T_134;
  wire [3:0] _T_136;
  wire [3:0] _T_138;
  wire [3:0] _T_140;
  wire  _T_145;
  wire [3:0] _T_146;
  wire  _T_147;
  wire [3:0] _T_148;
  wire  _T_149;
  wire [4:0] _T_150;
  wire  _T_151;
  wire [4:0] _T_152;
  wire  _T_157;
  wire  _T_158;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire [2:0] _T_178_opcode;
  assign io_tl_in_0_a_ready = _T_88;
  assign io_tl_in_0_d_valid = _T_158;
  assign io_tl_in_0_d_bits_opcode = _T_178_opcode;
  assign io_tl_in_0_d_bits_param = 2'h0;
  assign io_tl_in_0_d_bits_size = acq_size;
  assign io_tl_in_0_d_bits_source = acq_source;
  assign io_tl_in_0_d_bits_sink = 1'h0;
  assign io_tl_in_0_d_bits_data = _GEN_4;
  assign io_tl_in_0_d_bits_error = 1'h0;
  assign io_dmem_req_valid = _T_87;
  assign io_dmem_req_bits_addr = _T_90_address;
  assign io_dmem_req_bits_tag = 7'h0;
  assign io_dmem_req_bits_cmd = _T_152;
  assign io_dmem_req_bits_typ = _T_92_typ;
  assign io_dmem_req_bits_phys = 1'h1;
  assign io_dmem_s1_kill = 1'h0;
  assign io_dmem_s1_data_data = acq_data;
  assign io_dmem_s1_data_mask = acq_mask;
  assign io_dmem_invalidate_lr = 1'h0;
  assign _GEN_0 = io_dmem_resp_valid ? 2'h3 : state;
  assign _T_80 = io_tl_in_0_d_ready & io_tl_in_0_d_valid;
  assign _GEN_1 = _T_80 ? 2'h0 : _GEN_0;
  assign _GEN_2 = io_dmem_s2_nack ? 2'h2 : _GEN_1;
  assign _T_81 = io_dmem_req_ready & io_dmem_req_valid;
  assign _GEN_3 = _T_81 ? 2'h1 : _GEN_2;
  assign _GEN_4 = io_dmem_resp_valid ? io_dmem_resp_bits_data_raw : acq_data;
  assign _T_82 = io_tl_in_0_a_ready & io_tl_in_0_a_valid;
  assign _GEN_5 = _T_82 ? io_tl_in_0_a_bits_opcode : acq_opcode;
  assign _GEN_6 = _T_82 ? io_tl_in_0_a_bits_param : acq_param;
  assign _GEN_7 = _T_82 ? io_tl_in_0_a_bits_size : acq_size;
  assign _GEN_8 = _T_82 ? io_tl_in_0_a_bits_source : acq_source;
  assign _GEN_9 = _T_82 ? io_tl_in_0_a_bits_address : acq_address;
  assign _GEN_10 = _T_82 ? io_tl_in_0_a_bits_mask : acq_mask;
  assign _GEN_11 = _T_82 ? io_tl_in_0_a_bits_data : _GEN_4;
  assign _T_83 = state == 2'h0;
  assign ready = _T_83 | _T_80;
  assign _T_85 = io_tl_in_0_a_valid & ready;
  assign _T_86 = state == 2'h2;
  assign _T_87 = _T_85 | _T_86;
  assign _T_88 = io_dmem_req_ready & ready;
  assign _T_90_opcode = _T_86 ? acq_opcode : io_tl_in_0_a_bits_opcode;
  assign _T_90_param = _T_86 ? acq_param : io_tl_in_0_a_bits_param;
  assign _T_90_size = _T_86 ? acq_size : io_tl_in_0_a_bits_size;
  assign _T_90_address = _T_86 ? acq_address : io_tl_in_0_a_bits_address;
  assign _T_92_typ = {{1'd0}, _T_90_size};
  assign _T_112 = 3'h4 == _T_90_param;
  assign _T_113 = _T_112 ? 4'h8 : 4'h0;
  assign _T_114 = 3'h3 == _T_90_param;
  assign _T_115 = _T_114 ? 4'hf : _T_113;
  assign _T_116 = 3'h2 == _T_90_param;
  assign _T_117 = _T_116 ? 4'he : _T_115;
  assign _T_118 = 3'h1 == _T_90_param;
  assign _T_119 = _T_118 ? 4'hd : _T_117;
  assign _T_120 = 3'h0 == _T_90_param;
  assign _T_121 = _T_120 ? 4'hc : _T_119;
  assign _T_134 = _T_114 ? 3'h4 : 3'h0;
  assign _T_136 = _T_116 ? 4'hb : {{1'd0}, _T_134};
  assign _T_138 = _T_118 ? 4'ha : _T_136;
  assign _T_140 = _T_120 ? 4'h9 : _T_138;
  assign _T_145 = 3'h3 == _T_90_opcode;
  assign _T_146 = _T_145 ? _T_140 : 4'h0;
  assign _T_147 = 3'h2 == _T_90_opcode;
  assign _T_148 = _T_147 ? _T_121 : _T_146;
  assign _T_149 = 3'h1 == _T_90_opcode;
  assign _T_150 = _T_149 ? 5'h11 : {{1'd0}, _T_148};
  assign _T_151 = 3'h0 == _T_90_opcode;
  assign _T_152 = _T_151 ? 5'h1 : _T_150;
  assign _T_157 = state == 2'h3;
  assign _T_158 = io_dmem_resp_valid | _T_157;
  assign _T_161 = acq_opcode == 3'h0;
  assign _T_162 = acq_opcode == 3'h1;
  assign _T_163 = _T_161 | _T_162;
  assign _T_178_opcode = _T_163 ? 3'h0 : 3'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  acq_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  acq_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  acq_size = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  acq_source = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  acq_address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  acq_mask = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  acq_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_81) begin
        state <= 2'h1;
      end else begin
        if (io_dmem_s2_nack) begin
          state <= 2'h2;
        end else begin
          if (_T_80) begin
            state <= 2'h0;
          end else begin
            if (io_dmem_resp_valid) begin
              state <= 2'h3;
            end
          end
        end
      end
    end
    if (_T_82) begin
      acq_opcode <= io_tl_in_0_a_bits_opcode;
    end
    if (_T_82) begin
      acq_param <= io_tl_in_0_a_bits_param;
    end
    if (_T_82) begin
      acq_size <= io_tl_in_0_a_bits_size;
    end
    if (_T_82) begin
      acq_source <= io_tl_in_0_a_bits_source;
    end
    if (_T_82) begin
      acq_address <= io_tl_in_0_a_bits_address;
    end
    if (_T_82) begin
      acq_mask <= io_tl_in_0_a_bits_mask;
    end
    if (_T_82) begin
      acq_data <= io_tl_in_0_a_bits_data;
    end else begin
      if (io_dmem_resp_valid) begin
        acq_data <= io_dmem_resp_bits_data_raw;
      end
    end
  end
endmodule
module Repeater_5(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_full,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [2:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [2:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] saved_param;
  reg [31:0] _RAND_2;
  reg [2:0] saved_size;
  reg [31:0] _RAND_3;
  reg [4:0] saved_source;
  reg [31:0] _RAND_4;
  reg [31:0] saved_address;
  reg [31:0] _RAND_5;
  reg [3:0] saved_mask;
  reg [31:0] _RAND_6;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [2:0] _T_20_param;
  wire [2:0] _T_20_size;
  wire [4:0] _T_20_source;
  wire [31:0] _T_20_address;
  wire [3:0] _T_20_mask;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_2;
  wire [2:0] _GEN_3;
  wire [4:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [3:0] _GEN_6;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_full = full;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_param = _T_20_param;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_address = _T_20_address;
  assign io_deq_bits_mask = _T_20_mask;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_param = full ? saved_param : io_enq_bits_param;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_address = full ? saved_address : io_enq_bits_address;
  assign _T_20_mask = full ? saved_mask : io_enq_bits_mask;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_2 = _T_22 ? io_enq_bits_param : saved_param;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_address : saved_address;
  assign _GEN_6 = _T_22 ? io_enq_bits_mask : saved_mask;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_size = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_source = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  saved_mask = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_22) begin
      saved_mask <= io_enq_bits_mask;
    end
  end
endmodule
module TLFragmenter_2(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [2:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [2:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [1:0]  io_out_0_a_bits_size,
  output [9:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [1:0]  io_out_0_d_bits_size,
  input  [9:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  reg [3:0] _T_92;
  reg [31:0] _RAND_0;
  reg [2:0] _T_94;
  reg [31:0] _RAND_1;
  reg  _T_97;
  reg [31:0] _RAND_2;
  wire [3:0] _T_98;
  wire  _T_100;
  wire [3:0] _T_105;
  wire [2:0] _T_106;
  wire [4:0] _T_109;
  wire [1:0] _T_110;
  wire [1:0] _T_111;
  wire  _T_112;
  wire  _T_116;
  wire  _T_128;
  wire  _T_129;
  wire [5:0] _GEN_7;
  wire [5:0] _T_130;
  wire [5:0] _GEN_8;
  wire [5:0] _T_131;
  wire [6:0] _GEN_9;
  wire [6:0] _T_132;
  wire [6:0] _T_134;
  wire [6:0] _T_136;
  wire [6:0] _T_137;
  wire [6:0] _T_138;
  wire [2:0] _T_139;
  wire [3:0] _T_140;
  wire  _T_142;
  wire [3:0] _GEN_10;
  wire [3:0] _T_143;
  wire [1:0] _T_144;
  wire [1:0] _T_145;
  wire  _T_147;
  wire [1:0] _T_148;
  wire  _T_149;
  wire [1:0] _T_150;
  wire [2:0] _T_151;
  wire  _T_152;
  wire [3:0] _GEN_11;
  wire [4:0] _T_153;
  wire [4:0] _T_154;
  wire [3:0] _T_155;
  wire [3:0] _T_156;
  wire  _T_157;
  wire [2:0] _GEN_0;
  wire  _GEN_1;
  wire [3:0] _GEN_2;
  wire [2:0] _GEN_3;
  wire  _GEN_4;
  wire  _T_159;
  wire  _T_161;
  wire  _T_162;
  wire  _T_163;
  wire  _T_165;
  wire  _T_166;
  wire [4:0] _T_167;
  wire  _T_172;
  wire  _T_173;
  wire  _T_176;
  wire  _T_177;
  wire  _T_179;
  wire  Repeater_clock;
  wire  Repeater_reset;
  wire  Repeater_io_repeat;
  wire  Repeater_io_full;
  wire  Repeater_io_enq_ready;
  wire  Repeater_io_enq_valid;
  wire [2:0] Repeater_io_enq_bits_opcode;
  wire [2:0] Repeater_io_enq_bits_param;
  wire [2:0] Repeater_io_enq_bits_size;
  wire [4:0] Repeater_io_enq_bits_source;
  wire [31:0] Repeater_io_enq_bits_address;
  wire [3:0] Repeater_io_enq_bits_mask;
  wire  Repeater_io_deq_ready;
  wire  Repeater_io_deq_valid;
  wire [2:0] Repeater_io_deq_bits_opcode;
  wire [2:0] Repeater_io_deq_bits_param;
  wire [2:0] Repeater_io_deq_bits_size;
  wire [4:0] Repeater_io_deq_bits_source;
  wire [31:0] Repeater_io_deq_bits_address;
  wire [3:0] Repeater_io_deq_bits_mask;
  wire  _T_218;
  wire [2:0] _T_219;
  wire [12:0] _T_222;
  wire [5:0] _T_223;
  wire [5:0] _T_224;
  wire [8:0] _T_227;
  wire [1:0] _T_228;
  wire [1:0] _T_229;
  wire  _T_230;
  wire  _T_232;
  reg [3:0] _T_237;
  reg [31:0] _RAND_3;
  wire  _T_239;
  wire [3:0] _T_240;
  wire [4:0] _T_242;
  wire [4:0] _T_243;
  wire [3:0] _T_244;
  wire [3:0] _T_245;
  wire [3:0] _T_246;
  wire [3:0] _T_249;
  reg  _T_258;
  reg [31:0] _RAND_4;
  wire  _GEN_5;
  wire  _T_261;
  wire  _T_262;
  wire [3:0] _GEN_6;
  wire  _T_264;
  wire  _T_266;
  wire  _T_267;
  wire [5:0] _GEN_12;
  wire [5:0] _T_268;
  wire [5:0] _T_269;
  wire [5:0] _T_270;
  wire [5:0] _GEN_13;
  wire [5:0] _T_271;
  wire [5:0] _T_273;
  wire [5:0] _T_274;
  wire [31:0] _GEN_14;
  wire [31:0] _T_275;
  wire [5:0] _T_276;
  wire [9:0] _T_277;
  wire  _T_279;
  wire  _T_282;
  wire  _T_283;
  wire  _T_285;
  wire  _T_289;
  wire  _T_290;
  wire  _T_291;
  wire  _T_293;
  wire [3:0] _T_294;
  Repeater_5 Repeater (
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_full(Repeater_io_full),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_io_enq_bits_param),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_address(Repeater_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_io_enq_bits_mask),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_io_deq_bits_param),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_address(Repeater_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_io_deq_bits_mask)
  );
  assign io_in_0_a_ready = Repeater_io_enq_ready;
  assign io_in_0_d_valid = _T_166;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_param = io_out_0_d_bits_param;
  assign io_in_0_d_bits_size = _GEN_0;
  assign io_in_0_d_bits_source = _T_167;
  assign io_in_0_d_bits_sink = io_out_0_d_bits_sink;
  assign io_in_0_d_bits_data = io_out_0_d_bits_data;
  assign io_in_0_d_bits_error = io_out_0_d_bits_error;
  assign io_out_0_a_valid = Repeater_io_deq_valid;
  assign io_out_0_a_bits_opcode = Repeater_io_deq_bits_opcode;
  assign io_out_0_a_bits_param = Repeater_io_deq_bits_param;
  assign io_out_0_a_bits_size = _T_219[1:0];
  assign io_out_0_a_bits_source = _T_277;
  assign io_out_0_a_bits_address = _T_275;
  assign io_out_0_a_bits_mask = _T_294;
  assign io_out_0_a_bits_data = io_in_0_a_bits_data;
  assign io_out_0_d_ready = _T_163;
  assign _T_98 = io_out_0_d_bits_source[3:0];
  assign _T_100 = _T_92 == 4'h0;
  assign _T_105 = 4'h1 << io_out_0_d_bits_size;
  assign _T_106 = _T_105[2:0];
  assign _T_109 = 5'h3 << io_out_0_d_bits_size;
  assign _T_110 = _T_109[1:0];
  assign _T_111 = ~ _T_110;
  assign _T_112 = io_out_0_d_bits_opcode[0];
  assign _T_116 = io_out_0_d_valid == 1'h0;
  assign _T_128 = _T_106[2:2];
  assign _T_129 = _T_112 ? 1'h1 : _T_128;
  assign _GEN_7 = {{2'd0}, _T_98};
  assign _T_130 = _GEN_7 << 2;
  assign _GEN_8 = {{4'd0}, _T_111};
  assign _T_131 = _T_130 | _GEN_8;
  assign _GEN_9 = {{1'd0}, _T_131};
  assign _T_132 = _GEN_9 << 1;
  assign _T_134 = _T_132 | 7'h1;
  assign _T_136 = {1'h0,_T_131};
  assign _T_137 = ~ _T_136;
  assign _T_138 = _T_134 & _T_137;
  assign _T_139 = _T_138[6:4];
  assign _T_140 = _T_138[3:0];
  assign _T_142 = _T_139 != 3'h0;
  assign _GEN_10 = {{1'd0}, _T_139};
  assign _T_143 = _GEN_10 | _T_140;
  assign _T_144 = _T_143[3:2];
  assign _T_145 = _T_143[1:0];
  assign _T_147 = _T_144 != 2'h0;
  assign _T_148 = _T_144 | _T_145;
  assign _T_149 = _T_148[1];
  assign _T_150 = {_T_147,_T_149};
  assign _T_151 = {_T_142,_T_150};
  assign _T_152 = io_out_0_d_ready & io_out_0_d_valid;
  assign _GEN_11 = {{3'd0}, _T_129};
  assign _T_153 = _T_92 - _GEN_11;
  assign _T_154 = $unsigned(_T_153);
  assign _T_155 = _T_154[3:0];
  assign _T_156 = _T_100 ? _T_98 : _T_155;
  assign _T_157 = io_out_0_d_bits_source[4];
  assign _GEN_0 = _T_100 ? _T_151 : _T_94;
  assign _GEN_1 = _T_100 ? _T_157 : _T_97;
  assign _GEN_2 = _T_152 ? _T_156 : _T_92;
  assign _GEN_3 = _T_152 ? _GEN_0 : _T_94;
  assign _GEN_4 = _T_152 ? _GEN_1 : _T_97;
  assign _T_159 = _T_112 == 1'h0;
  assign _T_161 = _T_100 == 1'h0;
  assign _T_162 = _T_159 & _T_161;
  assign _T_163 = io_in_0_d_ready | _T_162;
  assign _T_165 = _T_162 == 1'h0;
  assign _T_166 = io_out_0_d_valid & _T_165;
  assign _T_167 = io_out_0_d_bits_source[9:5];
  assign _T_172 = io_out_0_d_bits_error == 1'h0;
  assign _T_173 = _T_116 | _T_172;
  assign _T_176 = _T_173 | _T_165;
  assign _T_177 = _T_176 | reset;
  assign _T_179 = _T_177 == 1'h0;
  assign Repeater_clock = clock;
  assign Repeater_reset = reset;
  assign Repeater_io_repeat = _T_267;
  assign Repeater_io_enq_valid = io_in_0_a_valid;
  assign Repeater_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Repeater_io_enq_bits_param = io_in_0_a_bits_param;
  assign Repeater_io_enq_bits_size = io_in_0_a_bits_size;
  assign Repeater_io_enq_bits_source = io_in_0_a_bits_source;
  assign Repeater_io_enq_bits_address = io_in_0_a_bits_address;
  assign Repeater_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Repeater_io_deq_ready = io_out_0_a_ready;
  assign _T_218 = Repeater_io_deq_bits_size > 3'h2;
  assign _T_219 = _T_218 ? 3'h2 : Repeater_io_deq_bits_size;
  assign _T_222 = 13'h3f << Repeater_io_deq_bits_size;
  assign _T_223 = _T_222[5:0];
  assign _T_224 = ~ _T_223;
  assign _T_227 = 9'h3 << _T_219;
  assign _T_228 = _T_227[1:0];
  assign _T_229 = ~ _T_228;
  assign _T_230 = Repeater_io_deq_bits_opcode[2];
  assign _T_232 = _T_230 == 1'h0;
  assign _T_239 = _T_237 == 4'h0;
  assign _T_240 = _T_224[5:2];
  assign _T_242 = _T_237 - 4'h1;
  assign _T_243 = $unsigned(_T_242);
  assign _T_244 = _T_243[3:0];
  assign _T_245 = _T_239 ? _T_240 : _T_244;
  assign _T_246 = ~ _T_245;
  assign _T_249 = ~ _T_246;
  assign _GEN_5 = _T_239 ? _T_97 : _T_258;
  assign _T_261 = _GEN_5 == 1'h0;
  assign _T_262 = io_out_0_a_ready & io_out_0_a_valid;
  assign _GEN_6 = _T_262 ? _T_249 : _T_237;
  assign _T_264 = _T_232 == 1'h0;
  assign _T_266 = _T_249 != 4'h0;
  assign _T_267 = _T_264 & _T_266;
  assign _GEN_12 = {{2'd0}, _T_245};
  assign _T_268 = _GEN_12 << 2;
  assign _T_269 = ~ _T_224;
  assign _T_270 = _T_268 | _T_269;
  assign _GEN_13 = {{4'd0}, _T_229};
  assign _T_271 = _T_270 | _GEN_13;
  assign _T_273 = _T_271 | 6'h3;
  assign _T_274 = ~ _T_273;
  assign _GEN_14 = {{26'd0}, _T_274};
  assign _T_275 = Repeater_io_deq_bits_address | _GEN_14;
  assign _T_276 = {Repeater_io_deq_bits_source,_T_261};
  assign _T_277 = {_T_276,_T_249};
  assign _T_279 = Repeater_io_full == 1'h0;
  assign _T_282 = _T_279 | _T_264;
  assign _T_283 = _T_282 | reset;
  assign _T_285 = _T_283 == 1'h0;
  assign _T_289 = Repeater_io_deq_bits_mask == 4'hf;
  assign _T_290 = _T_279 | _T_289;
  assign _T_291 = _T_290 | reset;
  assign _T_293 = _T_291 == 1'h0;
  assign _T_294 = Repeater_io_full ? 4'hf : io_in_0_a_bits_mask;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_92 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_94 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_97 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_237 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_258 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_92 <= 4'h0;
    end else begin
      if (_T_152) begin
        if (_T_100) begin
          _T_92 <= _T_98;
        end else begin
          _T_92 <= _T_155;
        end
      end
    end
    if (_T_152) begin
      if (_T_100) begin
        _T_94 <= _T_151;
      end
    end
    if (reset) begin
      _T_97 <= 1'h0;
    end else begin
      if (_T_152) begin
        if (_T_100) begin
          _T_97 <= _T_157;
        end
      end
    end
    if (reset) begin
      _T_237 <= 4'h0;
    end else begin
      if (_T_262) begin
        _T_237 <= _T_249;
      end
    end
    if (_T_239) begin
      _T_258 <= _T_97;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:174 assert (!out.d.valid || (acknum_fragment & acknum_size) === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_179) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:199 assert (!out.d.valid || !out.d.bits.error || !drop)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_285) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:273 assert (!repeater.io.full || !aHasData)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_285) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_293) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:276 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_293) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module HellaCacheArbiter(
  input         clock,
  output        io_requestor_0_req_ready,
  input         io_requestor_0_req_valid,
  input  [31:0] io_requestor_0_req_bits_addr,
  input  [6:0]  io_requestor_0_req_bits_tag,
  input  [4:0]  io_requestor_0_req_bits_cmd,
  input  [2:0]  io_requestor_0_req_bits_typ,
  input         io_requestor_0_req_bits_phys,
  input         io_requestor_0_s1_kill,
  input  [31:0] io_requestor_0_s1_data_data,
  input  [3:0]  io_requestor_0_s1_data_mask,
  output        io_requestor_0_s2_nack,
  output        io_requestor_0_resp_valid,
  output [31:0] io_requestor_0_resp_bits_data_raw,
  input         io_requestor_0_invalidate_lr,
  output        io_requestor_1_req_ready,
  input         io_requestor_1_req_valid,
  input  [31:0] io_requestor_1_req_bits_addr,
  input  [6:0]  io_requestor_1_req_bits_tag,
  input  [4:0]  io_requestor_1_req_bits_cmd,
  input  [2:0]  io_requestor_1_req_bits_typ,
  input         io_requestor_1_req_bits_phys,
  input         io_requestor_1_s1_kill,
  input  [31:0] io_requestor_1_s1_data_data,
  input  [3:0]  io_requestor_1_s1_data_mask,
  output        io_requestor_1_s2_nack,
  output        io_requestor_1_resp_valid,
  output [6:0]  io_requestor_1_resp_bits_tag,
  output [31:0] io_requestor_1_resp_bits_data,
  output        io_requestor_1_resp_bits_replay,
  output        io_requestor_1_resp_bits_has_data,
  output [31:0] io_requestor_1_resp_bits_data_word_bypass,
  output        io_requestor_1_replay_next,
  output        io_requestor_1_s2_xcpt_ma_ld,
  output        io_requestor_1_s2_xcpt_ma_st,
  output        io_requestor_1_s2_xcpt_pf_ld,
  output        io_requestor_1_s2_xcpt_pf_st,
  output        io_requestor_1_s2_xcpt_ae_ld,
  output        io_requestor_1_s2_xcpt_ae_st,
  input         io_requestor_1_invalidate_lr,
  output        io_requestor_1_ordered,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [6:0]  io_mem_req_bits_tag,
  output [4:0]  io_mem_req_bits_cmd,
  output [2:0]  io_mem_req_bits_typ,
  output        io_mem_req_bits_phys,
  output        io_mem_s1_kill,
  output [31:0] io_mem_s1_data_data,
  output [3:0]  io_mem_s1_data_mask,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [6:0]  io_mem_resp_bits_tag,
  input  [31:0] io_mem_resp_bits_data,
  input         io_mem_resp_bits_replay,
  input         io_mem_resp_bits_has_data,
  input  [31:0] io_mem_resp_bits_data_word_bypass,
  input  [31:0] io_mem_resp_bits_data_raw,
  input         io_mem_replay_next,
  input         io_mem_s2_xcpt_ma_ld,
  input         io_mem_s2_xcpt_ma_st,
  input         io_mem_s2_xcpt_pf_ld,
  input         io_mem_s2_xcpt_pf_st,
  input         io_mem_s2_xcpt_ae_ld,
  input         io_mem_s2_xcpt_ae_st,
  output        io_mem_invalidate_lr,
  input         io_mem_ordered
);
  reg  _T_208;
  reg [31:0] _RAND_0;
  reg  _T_210;
  reg [31:0] _RAND_1;
  wire  _T_211;
  wire  _T_212;
  wire  _T_214;
  wire  _T_215;
  wire [7:0] _T_217;
  wire [7:0] _T_220;
  wire [4:0] _GEN_0;
  wire [2:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire  _GEN_3;
  wire [7:0] _GEN_4;
  wire  _GEN_5;
  wire  _T_223;
  wire  _GEN_6;
  wire [31:0] _GEN_7;
  wire [3:0] _GEN_8;
  wire  _T_224;
  wire  _T_226;
  wire  _T_227;
  wire  _T_229;
  wire  _T_230;
  wire [5:0] _T_231;
  wire  _T_235;
  wire  _T_238;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_0_s2_nack = _T_230;
  assign io_requestor_0_resp_valid = _T_227;
  assign io_requestor_0_resp_bits_data_raw = io_mem_resp_bits_data_raw;
  assign io_requestor_1_req_ready = _T_215;
  assign io_requestor_1_s2_nack = _T_238;
  assign io_requestor_1_resp_valid = _T_235;
  assign io_requestor_1_resp_bits_tag = {{1'd0}, _T_231};
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_replay_next = io_mem_replay_next;
  assign io_requestor_1_s2_xcpt_ma_ld = io_mem_s2_xcpt_ma_ld;
  assign io_requestor_1_s2_xcpt_ma_st = io_mem_s2_xcpt_ma_st;
  assign io_requestor_1_s2_xcpt_pf_ld = io_mem_s2_xcpt_pf_ld;
  assign io_requestor_1_s2_xcpt_pf_st = io_mem_s2_xcpt_pf_st;
  assign io_requestor_1_s2_xcpt_ae_ld = io_mem_s2_xcpt_ae_ld;
  assign io_requestor_1_s2_xcpt_ae_st = io_mem_s2_xcpt_ae_st;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_mem_req_valid = _T_212;
  assign io_mem_req_bits_addr = _GEN_2;
  assign io_mem_req_bits_tag = _GEN_4[6:0];
  assign io_mem_req_bits_cmd = _GEN_0;
  assign io_mem_req_bits_typ = _GEN_1;
  assign io_mem_req_bits_phys = _GEN_3;
  assign io_mem_s1_kill = _GEN_6;
  assign io_mem_s1_data_data = _GEN_7;
  assign io_mem_s1_data_mask = _GEN_8;
  assign io_mem_invalidate_lr = _T_211;
  assign _T_211 = io_requestor_0_invalidate_lr | io_requestor_1_invalidate_lr;
  assign _T_212 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign _T_214 = io_requestor_0_req_valid == 1'h0;
  assign _T_215 = io_requestor_0_req_ready & _T_214;
  assign _T_217 = {io_requestor_1_req_bits_tag,1'h1};
  assign _T_220 = {io_requestor_0_req_bits_tag,1'h0};
  assign _GEN_0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign _GEN_1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign _GEN_2 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign _GEN_3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign _GEN_4 = io_requestor_0_req_valid ? _T_220 : _T_217;
  assign _GEN_5 = io_requestor_0_req_valid ? 1'h0 : 1'h1;
  assign _T_223 = _T_208 == 1'h0;
  assign _GEN_6 = _T_223 ? io_requestor_0_s1_kill : io_requestor_1_s1_kill;
  assign _GEN_7 = _T_223 ? io_requestor_0_s1_data_data : io_requestor_1_s1_data_data;
  assign _GEN_8 = _T_223 ? io_requestor_0_s1_data_mask : io_requestor_1_s1_data_mask;
  assign _T_224 = io_mem_resp_bits_tag[0];
  assign _T_226 = _T_224 == 1'h0;
  assign _T_227 = io_mem_resp_valid & _T_226;
  assign _T_229 = _T_210 == 1'h0;
  assign _T_230 = io_mem_s2_nack & _T_229;
  assign _T_231 = io_mem_resp_bits_tag[6:1];
  assign _T_235 = io_mem_resp_valid & _T_224;
  assign _T_238 = io_mem_s2_nack & _T_210;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_208 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_210 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_requestor_0_req_valid) begin
      _T_208 <= 1'h0;
    end else begin
      _T_208 <= 1'h1;
    end
    _T_210 <= _T_208;
  end
endmodule
module RRArbiter(
  input         clock,
  input         io_in_0_valid,
  input  [19:0] io_in_0_bits_addr,
  input         io_in_1_valid,
  input  [19:0] io_in_1_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [19:0] io_out_bits_addr,
  output        io_chosen
);
  wire  _GEN_3;
  wire [19:0] _GEN_4;
  wire  _T_60;
  reg  lastGrant;
  reg [31:0] _RAND_0;
  wire  _GEN_5;
  wire  grantMask_1;
  wire  validMask_1;
  wire  _GEN_6;
  wire  _GEN_7;
  assign io_out_valid = _GEN_3;
  assign io_out_bits_addr = _GEN_4;
  assign io_chosen = _GEN_7;
  assign _GEN_3 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign _GEN_4 = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign _T_60 = io_out_ready & io_out_valid;
  assign _GEN_5 = _T_60 ? io_chosen : lastGrant;
  assign grantMask_1 = 1'h1 > lastGrant;
  assign validMask_1 = io_in_1_valid & grantMask_1;
  assign _GEN_6 = io_in_0_valid ? 1'h0 : 1'h1;
  assign _GEN_7 = validMask_1 ? 1'h1 : _GEN_6;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  lastGrant = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_60) begin
      lastGrant <= io_chosen;
    end
  end
endmodule
module PTW(
  input         clock,
  input         reset,
  input         io_requestor_0_req_valid,
  input  [19:0] io_requestor_0_req_bits_addr,
  output        io_requestor_0_resp_valid,
  output [1:0]  io_requestor_0_status_dprv,
  output [1:0]  io_requestor_0_status_prv,
  output        io_requestor_0_status_mxr,
  output        io_requestor_0_status_sum,
  output        io_requestor_0_pmp_0_cfg_l,
  output [1:0]  io_requestor_0_pmp_0_cfg_a,
  output        io_requestor_0_pmp_0_cfg_x,
  output        io_requestor_0_pmp_0_cfg_w,
  output        io_requestor_0_pmp_0_cfg_r,
  output [29:0] io_requestor_0_pmp_0_addr,
  output [31:0] io_requestor_0_pmp_0_mask,
  output        io_requestor_0_pmp_1_cfg_l,
  output [1:0]  io_requestor_0_pmp_1_cfg_a,
  output        io_requestor_0_pmp_1_cfg_x,
  output        io_requestor_0_pmp_1_cfg_w,
  output        io_requestor_0_pmp_1_cfg_r,
  output [29:0] io_requestor_0_pmp_1_addr,
  output [31:0] io_requestor_0_pmp_1_mask,
  output        io_requestor_0_pmp_2_cfg_l,
  output [1:0]  io_requestor_0_pmp_2_cfg_a,
  output        io_requestor_0_pmp_2_cfg_x,
  output        io_requestor_0_pmp_2_cfg_w,
  output        io_requestor_0_pmp_2_cfg_r,
  output [29:0] io_requestor_0_pmp_2_addr,
  output [31:0] io_requestor_0_pmp_2_mask,
  output        io_requestor_0_pmp_3_cfg_l,
  output [1:0]  io_requestor_0_pmp_3_cfg_a,
  output        io_requestor_0_pmp_3_cfg_x,
  output        io_requestor_0_pmp_3_cfg_w,
  output        io_requestor_0_pmp_3_cfg_r,
  output [29:0] io_requestor_0_pmp_3_addr,
  output [31:0] io_requestor_0_pmp_3_mask,
  output        io_requestor_0_pmp_4_cfg_l,
  output [1:0]  io_requestor_0_pmp_4_cfg_a,
  output        io_requestor_0_pmp_4_cfg_x,
  output        io_requestor_0_pmp_4_cfg_w,
  output        io_requestor_0_pmp_4_cfg_r,
  output [29:0] io_requestor_0_pmp_4_addr,
  output [31:0] io_requestor_0_pmp_4_mask,
  output        io_requestor_0_pmp_5_cfg_l,
  output [1:0]  io_requestor_0_pmp_5_cfg_a,
  output        io_requestor_0_pmp_5_cfg_x,
  output        io_requestor_0_pmp_5_cfg_w,
  output        io_requestor_0_pmp_5_cfg_r,
  output [29:0] io_requestor_0_pmp_5_addr,
  output [31:0] io_requestor_0_pmp_5_mask,
  output        io_requestor_0_pmp_6_cfg_l,
  output [1:0]  io_requestor_0_pmp_6_cfg_a,
  output        io_requestor_0_pmp_6_cfg_x,
  output        io_requestor_0_pmp_6_cfg_w,
  output        io_requestor_0_pmp_6_cfg_r,
  output [29:0] io_requestor_0_pmp_6_addr,
  output [31:0] io_requestor_0_pmp_6_mask,
  output        io_requestor_0_pmp_7_cfg_l,
  output [1:0]  io_requestor_0_pmp_7_cfg_a,
  output        io_requestor_0_pmp_7_cfg_x,
  output        io_requestor_0_pmp_7_cfg_w,
  output        io_requestor_0_pmp_7_cfg_r,
  output [29:0] io_requestor_0_pmp_7_addr,
  output [31:0] io_requestor_0_pmp_7_mask,
  input         io_requestor_1_req_valid,
  input  [19:0] io_requestor_1_req_bits_addr,
  output        io_requestor_1_resp_valid,
  output [1:0]  io_requestor_1_status_dprv,
  output [1:0]  io_requestor_1_status_prv,
  output        io_requestor_1_status_mxr,
  output        io_requestor_1_status_sum,
  output        io_requestor_1_pmp_0_cfg_l,
  output [1:0]  io_requestor_1_pmp_0_cfg_a,
  output        io_requestor_1_pmp_0_cfg_x,
  output        io_requestor_1_pmp_0_cfg_w,
  output        io_requestor_1_pmp_0_cfg_r,
  output [29:0] io_requestor_1_pmp_0_addr,
  output [31:0] io_requestor_1_pmp_0_mask,
  output        io_requestor_1_pmp_1_cfg_l,
  output [1:0]  io_requestor_1_pmp_1_cfg_a,
  output        io_requestor_1_pmp_1_cfg_x,
  output        io_requestor_1_pmp_1_cfg_w,
  output        io_requestor_1_pmp_1_cfg_r,
  output [29:0] io_requestor_1_pmp_1_addr,
  output [31:0] io_requestor_1_pmp_1_mask,
  output        io_requestor_1_pmp_2_cfg_l,
  output [1:0]  io_requestor_1_pmp_2_cfg_a,
  output        io_requestor_1_pmp_2_cfg_x,
  output        io_requestor_1_pmp_2_cfg_w,
  output        io_requestor_1_pmp_2_cfg_r,
  output [29:0] io_requestor_1_pmp_2_addr,
  output [31:0] io_requestor_1_pmp_2_mask,
  output        io_requestor_1_pmp_3_cfg_l,
  output [1:0]  io_requestor_1_pmp_3_cfg_a,
  output        io_requestor_1_pmp_3_cfg_x,
  output        io_requestor_1_pmp_3_cfg_w,
  output        io_requestor_1_pmp_3_cfg_r,
  output [29:0] io_requestor_1_pmp_3_addr,
  output [31:0] io_requestor_1_pmp_3_mask,
  output        io_requestor_1_pmp_4_cfg_l,
  output [1:0]  io_requestor_1_pmp_4_cfg_a,
  output        io_requestor_1_pmp_4_cfg_x,
  output        io_requestor_1_pmp_4_cfg_w,
  output        io_requestor_1_pmp_4_cfg_r,
  output [29:0] io_requestor_1_pmp_4_addr,
  output [31:0] io_requestor_1_pmp_4_mask,
  output        io_requestor_1_pmp_5_cfg_l,
  output [1:0]  io_requestor_1_pmp_5_cfg_a,
  output        io_requestor_1_pmp_5_cfg_x,
  output        io_requestor_1_pmp_5_cfg_w,
  output        io_requestor_1_pmp_5_cfg_r,
  output [29:0] io_requestor_1_pmp_5_addr,
  output [31:0] io_requestor_1_pmp_5_mask,
  output        io_requestor_1_pmp_6_cfg_l,
  output [1:0]  io_requestor_1_pmp_6_cfg_a,
  output        io_requestor_1_pmp_6_cfg_x,
  output        io_requestor_1_pmp_6_cfg_w,
  output        io_requestor_1_pmp_6_cfg_r,
  output [29:0] io_requestor_1_pmp_6_addr,
  output [31:0] io_requestor_1_pmp_6_mask,
  output        io_requestor_1_pmp_7_cfg_l,
  output [1:0]  io_requestor_1_pmp_7_cfg_a,
  output        io_requestor_1_pmp_7_cfg_x,
  output        io_requestor_1_pmp_7_cfg_w,
  output        io_requestor_1_pmp_7_cfg_r,
  output [29:0] io_requestor_1_pmp_7_addr,
  output [31:0] io_requestor_1_pmp_7_mask,
  input         io_mem_req_ready,
  input         io_mem_s2_nack,
  input         io_mem_resp_valid,
  input  [31:0] io_mem_resp_bits_data,
  input         io_mem_s2_xcpt_ae_ld,
  input  [21:0] io_dpath_ptbr_ppn,
  input         io_dpath_sfence_valid,
  input         io_dpath_sfence_bits_rs1,
  input  [1:0]  io_dpath_status_dprv,
  input  [1:0]  io_dpath_status_prv,
  input         io_dpath_status_mxr,
  input         io_dpath_status_sum,
  input         io_dpath_pmp_0_cfg_l,
  input  [1:0]  io_dpath_pmp_0_cfg_a,
  input         io_dpath_pmp_0_cfg_x,
  input         io_dpath_pmp_0_cfg_w,
  input         io_dpath_pmp_0_cfg_r,
  input  [29:0] io_dpath_pmp_0_addr,
  input  [31:0] io_dpath_pmp_0_mask,
  input         io_dpath_pmp_1_cfg_l,
  input  [1:0]  io_dpath_pmp_1_cfg_a,
  input         io_dpath_pmp_1_cfg_x,
  input         io_dpath_pmp_1_cfg_w,
  input         io_dpath_pmp_1_cfg_r,
  input  [29:0] io_dpath_pmp_1_addr,
  input  [31:0] io_dpath_pmp_1_mask,
  input         io_dpath_pmp_2_cfg_l,
  input  [1:0]  io_dpath_pmp_2_cfg_a,
  input         io_dpath_pmp_2_cfg_x,
  input         io_dpath_pmp_2_cfg_w,
  input         io_dpath_pmp_2_cfg_r,
  input  [29:0] io_dpath_pmp_2_addr,
  input  [31:0] io_dpath_pmp_2_mask,
  input         io_dpath_pmp_3_cfg_l,
  input  [1:0]  io_dpath_pmp_3_cfg_a,
  input         io_dpath_pmp_3_cfg_x,
  input         io_dpath_pmp_3_cfg_w,
  input         io_dpath_pmp_3_cfg_r,
  input  [29:0] io_dpath_pmp_3_addr,
  input  [31:0] io_dpath_pmp_3_mask,
  input         io_dpath_pmp_4_cfg_l,
  input  [1:0]  io_dpath_pmp_4_cfg_a,
  input         io_dpath_pmp_4_cfg_x,
  input         io_dpath_pmp_4_cfg_w,
  input         io_dpath_pmp_4_cfg_r,
  input  [29:0] io_dpath_pmp_4_addr,
  input  [31:0] io_dpath_pmp_4_mask,
  input         io_dpath_pmp_5_cfg_l,
  input  [1:0]  io_dpath_pmp_5_cfg_a,
  input         io_dpath_pmp_5_cfg_x,
  input         io_dpath_pmp_5_cfg_w,
  input         io_dpath_pmp_5_cfg_r,
  input  [29:0] io_dpath_pmp_5_addr,
  input  [31:0] io_dpath_pmp_5_mask,
  input         io_dpath_pmp_6_cfg_l,
  input  [1:0]  io_dpath_pmp_6_cfg_a,
  input         io_dpath_pmp_6_cfg_x,
  input         io_dpath_pmp_6_cfg_w,
  input         io_dpath_pmp_6_cfg_r,
  input  [29:0] io_dpath_pmp_6_addr,
  input  [31:0] io_dpath_pmp_6_mask,
  input         io_dpath_pmp_7_cfg_l,
  input  [1:0]  io_dpath_pmp_7_cfg_a,
  input         io_dpath_pmp_7_cfg_x,
  input         io_dpath_pmp_7_cfg_w,
  input         io_dpath_pmp_7_cfg_r,
  input  [29:0] io_dpath_pmp_7_addr,
  input  [31:0] io_dpath_pmp_7_mask
);
  reg [1:0] state;
  reg [31:0] _RAND_0;
  reg  count;
  reg [31:0] _RAND_1;
  reg  resp_valid_0;
  reg [31:0] _RAND_2;
  reg  resp_valid_1;
  reg [31:0] _RAND_3;
  reg [19:0] r_req_addr;
  reg [31:0] _RAND_4;
  reg  r_req_dest;
  reg [31:0] _RAND_5;
  reg [53:0] r_pte_ppn;
  reg [63:0] _RAND_6;
  wire [9:0] _T_335;
  wire [9:0] vpn_idxs_1;
  wire [9:0] vpn_idx;
  wire  arb_clock;
  wire  arb_io_in_0_valid;
  wire [19:0] arb_io_in_0_bits_addr;
  wire  arb_io_in_1_valid;
  wire [19:0] arb_io_in_1_bits_addr;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [19:0] arb_io_out_bits_addr;
  wire  arb_io_chosen;
  wire  _T_340;
  wire [63:0] _T_345;
  wire  _T_347;
  wire  _T_348;
  wire  _T_349;
  wire [53:0] _T_355;
  wire [63:0] _T_360;
  wire  _T_361;
  wire  _T_362;
  wire  _T_363;
  wire  _T_364;
  wire [53:0] pte_ppn;
  wire [19:0] _T_372;
  wire  _T_373;
  wire  _T_374;
  wire  _T_376;
  wire [9:0] _T_377;
  wire  _T_379;
  wire  _T_380;
  wire  _GEN_5;
  wire  _GEN_6;
  wire [33:0] _T_382;
  wire  invalid_paddr;
  wire  _T_385;
  wire  _T_386;
  wire  _T_388;
  wire  _T_389;
  wire  _T_391;
  wire  _T_392;
  wire  _T_394;
  wire  _T_395;
  wire  _T_397;
  wire  traverse;
  wire [63:0] _T_398;
  wire [65:0] _GEN_106;
  wire [65:0] pte_addr;
  wire  _T_399;
  wire [19:0] _GEN_7;
  wire  _GEN_8;
  wire [53:0] _GEN_9;
  reg [3:0] _T_401;
  reg [31:0] _RAND_7;
  reg [3:0] _T_404;
  reg [31:0] _RAND_8;
  reg [31:0] _T_408_0;
  reg [31:0] _RAND_9;
  reg [31:0] _T_408_1;
  reg [31:0] _RAND_10;
  reg [31:0] _T_408_2;
  reg [31:0] _RAND_11;
  reg [31:0] _T_408_3;
  reg [31:0] _RAND_12;
  reg [19:0] _T_418_0;
  reg [31:0] _RAND_13;
  reg [19:0] _T_418_1;
  reg [31:0] _RAND_14;
  reg [19:0] _T_418_2;
  reg [31:0] _RAND_15;
  reg [19:0] _T_418_3;
  reg [31:0] _RAND_16;
  wire [65:0] _GEN_107;
  wire  _T_425;
  wire [65:0] _GEN_108;
  wire  _T_426;
  wire [65:0] _GEN_109;
  wire  _T_427;
  wire [65:0] _GEN_110;
  wire  _T_428;
  wire [1:0] _T_429;
  wire [1:0] _T_430;
  wire [3:0] _T_431;
  wire [3:0] _T_432;
  wire  _T_434;
  wire  _T_435;
  wire  _T_437;
  wire  _T_438;
  wire [3:0] _T_439;
  wire  _T_441;
  wire [3:0] _T_443;
  wire  _T_444;
  wire [1:0] _T_445;
  wire [3:0] _T_446;
  wire  _T_447;
  wire [2:0] _T_448;
  wire [1:0] _T_449;
  wire  _T_451;
  wire  _T_452;
  wire  _T_453;
  wire [1:0] _T_459;
  wire [1:0] _T_460;
  wire [1:0] _T_461;
  wire [1:0] _T_462;
  wire [3:0] _T_464;
  wire [3:0] _T_465;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_12;
  wire [31:0] _GEN_13;
  wire [19:0] _GEN_1;
  wire [19:0] _GEN_14;
  wire [19:0] _GEN_15;
  wire [19:0] _GEN_16;
  wire [19:0] _GEN_17;
  wire [3:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire [31:0] _GEN_21;
  wire [31:0] _GEN_22;
  wire [19:0] _GEN_23;
  wire [19:0] _GEN_24;
  wire [19:0] _GEN_25;
  wire [19:0] _GEN_26;
  wire  _T_468;
  wire  _T_469;
  wire [1:0] _T_470;
  wire [1:0] _T_471;
  wire  _T_473;
  wire [1:0] _T_474;
  wire  _T_475;
  wire [1:0] _T_476;
  wire  _T_478;
  wire  _T_480;
  wire [1:0] _T_482;
  wire [3:0] _GEN_111;
  wire [3:0] _T_483;
  wire [3:0] _T_484;
  wire [3:0] _T_485;
  wire [3:0] _T_486;
  wire [3:0] _T_487;
  wire [1:0] _T_488;
  wire  _T_489;
  wire  _T_491;
  wire [3:0] _T_493;
  wire [3:0] _T_494;
  wire [3:0] _T_495;
  wire [3:0] _T_496;
  wire [3:0] _T_497;
  wire [3:0] _T_498;
  wire [3:0] _GEN_27;
  wire  _T_501;
  wire  _T_502;
  wire [3:0] _GEN_28;
  wire  pte_cache_hit;
  wire  _T_506;
  wire  _T_507;
  wire  _T_508;
  wire  _T_509;
  wire [19:0] _T_512;
  wire [19:0] _T_514;
  wire [19:0] _T_516;
  wire [19:0] _T_518;
  wire [19:0] _T_519;
  wire [19:0] _T_520;
  wire [19:0] _T_521;
  wire  _T_1183;
  wire [1:0] _GEN_29;
  wire [1:0] _GEN_30;
  wire  _GEN_31;
  wire  _T_1186;
  wire [1:0] _T_1189;
  wire  _T_1190;
  wire  _GEN_33;
  wire [53:0] _GEN_34;
  wire  _T_1192;
  wire  _T_1193;
  wire [1:0] _GEN_35;
  wire  _GEN_37;
  wire [53:0] _GEN_38;
  wire [1:0] _GEN_39;
  wire  _T_1194;
  wire [1:0] _GEN_40;
  wire  _T_1195;
  wire [1:0] _GEN_41;
  wire [1:0] _GEN_42;
  wire  _GEN_43;
  wire  _T_1200;
  wire  _GEN_44;
  wire [1:0] _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire [53:0] _GEN_51;
  wire [1:0] _GEN_61;
  wire  _GEN_62;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _GEN_68;
  wire [1:0] _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire [1:0] _GEN_73;
  wire [53:0] _GEN_74;
  wire  _GEN_84;
  wire  _GEN_87;
  wire  _GEN_88;
  RRArbiter arb (
    .clock(arb_clock),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_chosen(arb_io_chosen)
  );
  assign io_requestor_0_resp_valid = resp_valid_0;
  assign io_requestor_0_status_dprv = io_dpath_status_dprv;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_mxr = io_dpath_status_mxr;
  assign io_requestor_0_status_sum = io_dpath_status_sum;
  assign io_requestor_0_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l;
  assign io_requestor_0_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a;
  assign io_requestor_0_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x;
  assign io_requestor_0_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w;
  assign io_requestor_0_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r;
  assign io_requestor_0_pmp_0_addr = io_dpath_pmp_0_addr;
  assign io_requestor_0_pmp_0_mask = io_dpath_pmp_0_mask;
  assign io_requestor_0_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l;
  assign io_requestor_0_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a;
  assign io_requestor_0_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x;
  assign io_requestor_0_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w;
  assign io_requestor_0_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r;
  assign io_requestor_0_pmp_1_addr = io_dpath_pmp_1_addr;
  assign io_requestor_0_pmp_1_mask = io_dpath_pmp_1_mask;
  assign io_requestor_0_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l;
  assign io_requestor_0_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a;
  assign io_requestor_0_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x;
  assign io_requestor_0_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w;
  assign io_requestor_0_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r;
  assign io_requestor_0_pmp_2_addr = io_dpath_pmp_2_addr;
  assign io_requestor_0_pmp_2_mask = io_dpath_pmp_2_mask;
  assign io_requestor_0_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l;
  assign io_requestor_0_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a;
  assign io_requestor_0_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x;
  assign io_requestor_0_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w;
  assign io_requestor_0_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r;
  assign io_requestor_0_pmp_3_addr = io_dpath_pmp_3_addr;
  assign io_requestor_0_pmp_3_mask = io_dpath_pmp_3_mask;
  assign io_requestor_0_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l;
  assign io_requestor_0_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a;
  assign io_requestor_0_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x;
  assign io_requestor_0_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w;
  assign io_requestor_0_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r;
  assign io_requestor_0_pmp_4_addr = io_dpath_pmp_4_addr;
  assign io_requestor_0_pmp_4_mask = io_dpath_pmp_4_mask;
  assign io_requestor_0_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l;
  assign io_requestor_0_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a;
  assign io_requestor_0_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x;
  assign io_requestor_0_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w;
  assign io_requestor_0_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r;
  assign io_requestor_0_pmp_5_addr = io_dpath_pmp_5_addr;
  assign io_requestor_0_pmp_5_mask = io_dpath_pmp_5_mask;
  assign io_requestor_0_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l;
  assign io_requestor_0_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a;
  assign io_requestor_0_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x;
  assign io_requestor_0_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w;
  assign io_requestor_0_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r;
  assign io_requestor_0_pmp_6_addr = io_dpath_pmp_6_addr;
  assign io_requestor_0_pmp_6_mask = io_dpath_pmp_6_mask;
  assign io_requestor_0_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l;
  assign io_requestor_0_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a;
  assign io_requestor_0_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x;
  assign io_requestor_0_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w;
  assign io_requestor_0_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r;
  assign io_requestor_0_pmp_7_addr = io_dpath_pmp_7_addr;
  assign io_requestor_0_pmp_7_mask = io_dpath_pmp_7_mask;
  assign io_requestor_1_resp_valid = resp_valid_1;
  assign io_requestor_1_status_dprv = io_dpath_status_dprv;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_mxr = io_dpath_status_mxr;
  assign io_requestor_1_status_sum = io_dpath_status_sum;
  assign io_requestor_1_pmp_0_cfg_l = io_dpath_pmp_0_cfg_l;
  assign io_requestor_1_pmp_0_cfg_a = io_dpath_pmp_0_cfg_a;
  assign io_requestor_1_pmp_0_cfg_x = io_dpath_pmp_0_cfg_x;
  assign io_requestor_1_pmp_0_cfg_w = io_dpath_pmp_0_cfg_w;
  assign io_requestor_1_pmp_0_cfg_r = io_dpath_pmp_0_cfg_r;
  assign io_requestor_1_pmp_0_addr = io_dpath_pmp_0_addr;
  assign io_requestor_1_pmp_0_mask = io_dpath_pmp_0_mask;
  assign io_requestor_1_pmp_1_cfg_l = io_dpath_pmp_1_cfg_l;
  assign io_requestor_1_pmp_1_cfg_a = io_dpath_pmp_1_cfg_a;
  assign io_requestor_1_pmp_1_cfg_x = io_dpath_pmp_1_cfg_x;
  assign io_requestor_1_pmp_1_cfg_w = io_dpath_pmp_1_cfg_w;
  assign io_requestor_1_pmp_1_cfg_r = io_dpath_pmp_1_cfg_r;
  assign io_requestor_1_pmp_1_addr = io_dpath_pmp_1_addr;
  assign io_requestor_1_pmp_1_mask = io_dpath_pmp_1_mask;
  assign io_requestor_1_pmp_2_cfg_l = io_dpath_pmp_2_cfg_l;
  assign io_requestor_1_pmp_2_cfg_a = io_dpath_pmp_2_cfg_a;
  assign io_requestor_1_pmp_2_cfg_x = io_dpath_pmp_2_cfg_x;
  assign io_requestor_1_pmp_2_cfg_w = io_dpath_pmp_2_cfg_w;
  assign io_requestor_1_pmp_2_cfg_r = io_dpath_pmp_2_cfg_r;
  assign io_requestor_1_pmp_2_addr = io_dpath_pmp_2_addr;
  assign io_requestor_1_pmp_2_mask = io_dpath_pmp_2_mask;
  assign io_requestor_1_pmp_3_cfg_l = io_dpath_pmp_3_cfg_l;
  assign io_requestor_1_pmp_3_cfg_a = io_dpath_pmp_3_cfg_a;
  assign io_requestor_1_pmp_3_cfg_x = io_dpath_pmp_3_cfg_x;
  assign io_requestor_1_pmp_3_cfg_w = io_dpath_pmp_3_cfg_w;
  assign io_requestor_1_pmp_3_cfg_r = io_dpath_pmp_3_cfg_r;
  assign io_requestor_1_pmp_3_addr = io_dpath_pmp_3_addr;
  assign io_requestor_1_pmp_3_mask = io_dpath_pmp_3_mask;
  assign io_requestor_1_pmp_4_cfg_l = io_dpath_pmp_4_cfg_l;
  assign io_requestor_1_pmp_4_cfg_a = io_dpath_pmp_4_cfg_a;
  assign io_requestor_1_pmp_4_cfg_x = io_dpath_pmp_4_cfg_x;
  assign io_requestor_1_pmp_4_cfg_w = io_dpath_pmp_4_cfg_w;
  assign io_requestor_1_pmp_4_cfg_r = io_dpath_pmp_4_cfg_r;
  assign io_requestor_1_pmp_4_addr = io_dpath_pmp_4_addr;
  assign io_requestor_1_pmp_4_mask = io_dpath_pmp_4_mask;
  assign io_requestor_1_pmp_5_cfg_l = io_dpath_pmp_5_cfg_l;
  assign io_requestor_1_pmp_5_cfg_a = io_dpath_pmp_5_cfg_a;
  assign io_requestor_1_pmp_5_cfg_x = io_dpath_pmp_5_cfg_x;
  assign io_requestor_1_pmp_5_cfg_w = io_dpath_pmp_5_cfg_w;
  assign io_requestor_1_pmp_5_cfg_r = io_dpath_pmp_5_cfg_r;
  assign io_requestor_1_pmp_5_addr = io_dpath_pmp_5_addr;
  assign io_requestor_1_pmp_5_mask = io_dpath_pmp_5_mask;
  assign io_requestor_1_pmp_6_cfg_l = io_dpath_pmp_6_cfg_l;
  assign io_requestor_1_pmp_6_cfg_a = io_dpath_pmp_6_cfg_a;
  assign io_requestor_1_pmp_6_cfg_x = io_dpath_pmp_6_cfg_x;
  assign io_requestor_1_pmp_6_cfg_w = io_dpath_pmp_6_cfg_w;
  assign io_requestor_1_pmp_6_cfg_r = io_dpath_pmp_6_cfg_r;
  assign io_requestor_1_pmp_6_addr = io_dpath_pmp_6_addr;
  assign io_requestor_1_pmp_6_mask = io_dpath_pmp_6_mask;
  assign io_requestor_1_pmp_7_cfg_l = io_dpath_pmp_7_cfg_l;
  assign io_requestor_1_pmp_7_cfg_a = io_dpath_pmp_7_cfg_a;
  assign io_requestor_1_pmp_7_cfg_x = io_dpath_pmp_7_cfg_x;
  assign io_requestor_1_pmp_7_cfg_w = io_dpath_pmp_7_cfg_w;
  assign io_requestor_1_pmp_7_cfg_r = io_dpath_pmp_7_cfg_r;
  assign io_requestor_1_pmp_7_addr = io_dpath_pmp_7_addr;
  assign io_requestor_1_pmp_7_mask = io_dpath_pmp_7_mask;
  assign _T_335 = r_req_addr[19:10];
  assign vpn_idxs_1 = r_req_addr[9:0];
  assign vpn_idx = count ? vpn_idxs_1 : _T_335;
  assign arb_clock = clock;
  assign arb_io_in_0_valid = io_requestor_0_req_valid;
  assign arb_io_in_0_bits_addr = io_requestor_0_req_bits_addr;
  assign arb_io_in_1_valid = io_requestor_1_req_valid;
  assign arb_io_in_1_bits_addr = io_requestor_1_req_bits_addr;
  assign arb_io_out_ready = _T_340;
  assign _T_340 = state == 2'h0;
  assign _T_345 = {{32'd0}, io_mem_resp_bits_data};
  assign _T_347 = _T_345[1];
  assign _T_348 = _T_345[2];
  assign _T_349 = _T_345[3];
  assign _T_355 = _T_345[63:10];
  assign _T_360 = {{32'd0}, io_mem_resp_bits_data};
  assign _T_361 = _T_360[0];
  assign _T_362 = _T_360[1];
  assign _T_363 = _T_360[2];
  assign _T_364 = _T_360[3];
  assign pte_ppn = {{34'd0}, _T_372};
  assign _T_372 = _T_355[19:0];
  assign _T_373 = _T_347 | _T_348;
  assign _T_374 = _T_373 | _T_349;
  assign _T_376 = count <= 1'h0;
  assign _T_377 = _T_355[9:0];
  assign _T_379 = _T_377 != 10'h0;
  assign _T_380 = _T_376 & _T_379;
  assign _GEN_5 = _T_380 ? 1'h0 : _T_361;
  assign _GEN_6 = _T_374 ? _GEN_5 : _T_361;
  assign _T_382 = _T_355[53:20];
  assign invalid_paddr = _T_382 != 34'h0;
  assign _T_385 = _T_362 == 1'h0;
  assign _T_386 = _GEN_6 & _T_385;
  assign _T_388 = _T_363 == 1'h0;
  assign _T_389 = _T_386 & _T_388;
  assign _T_391 = _T_364 == 1'h0;
  assign _T_392 = _T_389 & _T_391;
  assign _T_394 = invalid_paddr == 1'h0;
  assign _T_395 = _T_392 & _T_394;
  assign _T_397 = count < 1'h1;
  assign traverse = _T_395 & _T_397;
  assign _T_398 = {r_pte_ppn,vpn_idx};
  assign _GEN_106 = {{2'd0}, _T_398};
  assign pte_addr = _GEN_106 << 2;
  assign _T_399 = arb_io_out_ready & arb_io_out_valid;
  assign _GEN_7 = _T_399 ? arb_io_out_bits_addr : r_req_addr;
  assign _GEN_8 = _T_399 ? arb_io_chosen : r_req_dest;
  assign _GEN_9 = _T_399 ? {{32'd0}, io_dpath_ptbr_ppn} : r_pte_ppn;
  assign _GEN_107 = {{34'd0}, _T_408_0};
  assign _T_425 = _GEN_107 == pte_addr;
  assign _GEN_108 = {{34'd0}, _T_408_1};
  assign _T_426 = _GEN_108 == pte_addr;
  assign _GEN_109 = {{34'd0}, _T_408_2};
  assign _T_427 = _GEN_109 == pte_addr;
  assign _GEN_110 = {{34'd0}, _T_408_3};
  assign _T_428 = _GEN_110 == pte_addr;
  assign _T_429 = {_T_426,_T_425};
  assign _T_430 = {_T_428,_T_427};
  assign _T_431 = {_T_430,_T_429};
  assign _T_432 = _T_431 & _T_404;
  assign _T_434 = _T_432 != 4'h0;
  assign _T_435 = io_mem_resp_valid & traverse;
  assign _T_437 = _T_434 == 1'h0;
  assign _T_438 = _T_435 & _T_437;
  assign _T_439 = ~ _T_404;
  assign _T_441 = _T_439 == 4'h0;
  assign _T_443 = _T_401 >> 1'h1;
  assign _T_444 = _T_443[0];
  assign _T_445 = {1'h1,_T_444};
  assign _T_446 = _T_401 >> _T_445;
  assign _T_447 = _T_446[0];
  assign _T_448 = {_T_445,_T_447};
  assign _T_449 = _T_448[1:0];
  assign _T_451 = _T_439[0];
  assign _T_452 = _T_439[1];
  assign _T_453 = _T_439[2];
  assign _T_459 = _T_453 ? 2'h2 : 2'h3;
  assign _T_460 = _T_452 ? 2'h1 : _T_459;
  assign _T_461 = _T_451 ? 2'h0 : _T_460;
  assign _T_462 = _T_441 ? _T_449 : _T_461;
  assign _T_464 = 4'h1 << _T_462;
  assign _T_465 = _T_404 | _T_464;
  assign _GEN_0 = pte_addr[31:0];
  assign _GEN_10 = 2'h0 == _T_462 ? _GEN_0 : _T_408_0;
  assign _GEN_11 = 2'h1 == _T_462 ? _GEN_0 : _T_408_1;
  assign _GEN_12 = 2'h2 == _T_462 ? _GEN_0 : _T_408_2;
  assign _GEN_13 = 2'h3 == _T_462 ? _GEN_0 : _T_408_3;
  assign _GEN_1 = pte_ppn[19:0];
  assign _GEN_14 = 2'h0 == _T_462 ? _GEN_1 : _T_418_0;
  assign _GEN_15 = 2'h1 == _T_462 ? _GEN_1 : _T_418_1;
  assign _GEN_16 = 2'h2 == _T_462 ? _GEN_1 : _T_418_2;
  assign _GEN_17 = 2'h3 == _T_462 ? _GEN_1 : _T_418_3;
  assign _GEN_18 = _T_438 ? _T_465 : _T_404;
  assign _GEN_19 = _T_438 ? _GEN_10 : _T_408_0;
  assign _GEN_20 = _T_438 ? _GEN_11 : _T_408_1;
  assign _GEN_21 = _T_438 ? _GEN_12 : _T_408_2;
  assign _GEN_22 = _T_438 ? _GEN_13 : _T_408_3;
  assign _GEN_23 = _T_438 ? _GEN_14 : _T_418_0;
  assign _GEN_24 = _T_438 ? _GEN_15 : _T_418_1;
  assign _GEN_25 = _T_438 ? _GEN_16 : _T_418_2;
  assign _GEN_26 = _T_438 ? _GEN_17 : _T_418_3;
  assign _T_468 = state == 2'h1;
  assign _T_469 = _T_434 & _T_468;
  assign _T_470 = _T_432[3:2];
  assign _T_471 = _T_432[1:0];
  assign _T_473 = _T_470 != 2'h0;
  assign _T_474 = _T_470 | _T_471;
  assign _T_475 = _T_474[1];
  assign _T_476 = {_T_473,_T_475};
  assign _T_478 = _T_476[1];
  assign _T_480 = _T_478 == 1'h0;
  assign _T_482 = 2'h1 << 1'h1;
  assign _GEN_111 = {{2'd0}, _T_482};
  assign _T_483 = _T_401 | _GEN_111;
  assign _T_484 = ~ _T_401;
  assign _T_485 = _T_484 | _GEN_111;
  assign _T_486 = ~ _T_485;
  assign _T_487 = _T_480 ? _T_483 : _T_486;
  assign _T_488 = {1'h1,_T_478};
  assign _T_489 = _T_476[0];
  assign _T_491 = _T_489 == 1'h0;
  assign _T_493 = 4'h1 << _T_488;
  assign _T_494 = _T_487 | _T_493;
  assign _T_495 = ~ _T_487;
  assign _T_496 = _T_495 | _T_493;
  assign _T_497 = ~ _T_496;
  assign _T_498 = _T_491 ? _T_494 : _T_497;
  assign _GEN_27 = _T_469 ? _T_498 : _T_401;
  assign _T_501 = io_dpath_sfence_bits_rs1 == 1'h0;
  assign _T_502 = io_dpath_sfence_valid & _T_501;
  assign _GEN_28 = _T_502 ? 4'h0 : _GEN_18;
  assign pte_cache_hit = _T_434 & _T_397;
  assign _T_506 = _T_432[0];
  assign _T_507 = _T_432[1];
  assign _T_508 = _T_432[2];
  assign _T_509 = _T_432[3];
  assign _T_512 = _T_506 ? _T_418_0 : 20'h0;
  assign _T_514 = _T_507 ? _T_418_1 : 20'h0;
  assign _T_516 = _T_508 ? _T_418_2 : 20'h0;
  assign _T_518 = _T_509 ? _T_418_3 : 20'h0;
  assign _T_519 = _T_512 | _T_514;
  assign _T_520 = _T_519 | _T_516;
  assign _T_521 = _T_520 | _T_518;
  assign _T_1183 = 2'h0 == state;
  assign _GEN_29 = _T_399 ? 2'h1 : state;
  assign _GEN_30 = _T_1183 ? _GEN_29 : state;
  assign _GEN_31 = _T_1183 ? 1'h0 : count;
  assign _T_1186 = 2'h1 == state;
  assign _T_1189 = count + 1'h1;
  assign _T_1190 = _T_1189[0:0];
  assign _GEN_33 = pte_cache_hit ? _T_1190 : _GEN_31;
  assign _GEN_34 = pte_cache_hit ? {{34'd0}, _T_521} : _GEN_9;
  assign _T_1192 = pte_cache_hit == 1'h0;
  assign _T_1193 = _T_1192 & io_mem_req_ready;
  assign _GEN_35 = _T_1193 ? 2'h2 : _GEN_30;
  assign _GEN_37 = _T_1186 ? _GEN_33 : _GEN_31;
  assign _GEN_38 = _T_1186 ? _GEN_34 : _GEN_9;
  assign _GEN_39 = _T_1186 ? _GEN_35 : _GEN_30;
  assign _T_1194 = 2'h2 == state;
  assign _GEN_40 = _T_1194 ? 2'h3 : _GEN_39;
  assign _T_1195 = 2'h3 == state;
  assign _GEN_41 = io_mem_s2_nack ? 2'h1 : _GEN_40;
  assign _GEN_42 = traverse ? 2'h1 : _GEN_41;
  assign _GEN_43 = traverse ? _T_1190 : _GEN_37;
  assign _T_1200 = traverse == 1'h0;
  assign _GEN_44 = 1'h0 == r_req_dest;
  assign _GEN_48 = _T_1200 ? 2'h0 : _GEN_42;
  assign _GEN_49 = _T_1200 ? _GEN_44 : 1'h0;
  assign _GEN_50 = _T_1200 ? r_req_dest : 1'h0;
  assign _GEN_51 = io_mem_resp_valid ? pte_ppn : _GEN_38;
  assign _GEN_61 = io_mem_resp_valid ? _GEN_48 : _GEN_41;
  assign _GEN_62 = io_mem_resp_valid ? _GEN_43 : _GEN_37;
  assign _GEN_65 = io_mem_resp_valid ? _GEN_49 : 1'h0;
  assign _GEN_66 = io_mem_resp_valid ? _GEN_50 : 1'h0;
  assign _GEN_67 = 1'h0 == r_req_dest ? 1'h1 : _GEN_65;
  assign _GEN_68 = r_req_dest ? 1'h1 : _GEN_66;
  assign _GEN_70 = io_mem_s2_xcpt_ae_ld ? 2'h0 : _GEN_61;
  assign _GEN_71 = io_mem_s2_xcpt_ae_ld ? _GEN_67 : _GEN_65;
  assign _GEN_72 = io_mem_s2_xcpt_ae_ld ? _GEN_68 : _GEN_66;
  assign _GEN_73 = _T_1195 ? _GEN_70 : _GEN_40;
  assign _GEN_74 = _T_1195 ? _GEN_51 : _GEN_38;
  assign _GEN_84 = _T_1195 ? _GEN_62 : _GEN_37;
  assign _GEN_87 = _T_1195 ? _GEN_71 : 1'h0;
  assign _GEN_88 = _T_1195 ? _GEN_72 : 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  count = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  resp_valid_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  resp_valid_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  r_req_addr = _RAND_4[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  r_req_dest = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{$random}};
  r_pte_ppn = _RAND_6[53:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_401 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_404 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_408_0 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_408_1 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_408_2 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_408_3 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_418_0 = _RAND_13[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_418_1 = _RAND_14[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_418_2 = _RAND_15[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_418_3 = _RAND_16[19:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_1195) begin
        if (io_mem_s2_xcpt_ae_ld) begin
          state <= 2'h0;
        end else begin
          if (io_mem_resp_valid) begin
            if (_T_1200) begin
              state <= 2'h0;
            end else begin
              if (traverse) begin
                state <= 2'h1;
              end else begin
                if (io_mem_s2_nack) begin
                  state <= 2'h1;
                end else begin
                  if (_T_1194) begin
                    state <= 2'h3;
                  end else begin
                    if (_T_1186) begin
                      if (_T_1193) begin
                        state <= 2'h2;
                      end else begin
                        if (_T_1183) begin
                          if (_T_399) begin
                            state <= 2'h1;
                          end
                        end
                      end
                    end else begin
                      if (_T_1183) begin
                        if (_T_399) begin
                          state <= 2'h1;
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (io_mem_s2_nack) begin
              state <= 2'h1;
            end else begin
              if (_T_1194) begin
                state <= 2'h3;
              end else begin
                if (_T_1186) begin
                  if (_T_1193) begin
                    state <= 2'h2;
                  end else begin
                    if (_T_1183) begin
                      if (_T_399) begin
                        state <= 2'h1;
                      end
                    end
                  end
                end else begin
                  if (_T_1183) begin
                    if (_T_399) begin
                      state <= 2'h1;
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_1194) begin
          state <= 2'h3;
        end else begin
          if (_T_1186) begin
            if (_T_1193) begin
              state <= 2'h2;
            end else begin
              state <= _GEN_30;
            end
          end else begin
            state <= _GEN_30;
          end
        end
      end
    end
    if (_T_1195) begin
      if (io_mem_resp_valid) begin
        if (traverse) begin
          count <= _T_1190;
        end else begin
          if (_T_1186) begin
            if (pte_cache_hit) begin
              count <= _T_1190;
            end else begin
              if (_T_1183) begin
                count <= 1'h0;
              end
            end
          end else begin
            if (_T_1183) begin
              count <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_1186) begin
          if (pte_cache_hit) begin
            count <= _T_1190;
          end else begin
            if (_T_1183) begin
              count <= 1'h0;
            end
          end
        end else begin
          if (_T_1183) begin
            count <= 1'h0;
          end
        end
      end
    end else begin
      if (_T_1186) begin
        if (pte_cache_hit) begin
          count <= _T_1190;
        end else begin
          count <= _GEN_31;
        end
      end else begin
        count <= _GEN_31;
      end
    end
    if (_T_1195) begin
      if (io_mem_s2_xcpt_ae_ld) begin
        if (1'h0 == r_req_dest) begin
          resp_valid_0 <= 1'h1;
        end else begin
          if (io_mem_resp_valid) begin
            if (_T_1200) begin
              resp_valid_0 <= _GEN_44;
            end else begin
              resp_valid_0 <= 1'h0;
            end
          end else begin
            resp_valid_0 <= 1'h0;
          end
        end
      end else begin
        if (io_mem_resp_valid) begin
          if (_T_1200) begin
            resp_valid_0 <= _GEN_44;
          end else begin
            resp_valid_0 <= 1'h0;
          end
        end else begin
          resp_valid_0 <= 1'h0;
        end
      end
    end else begin
      resp_valid_0 <= 1'h0;
    end
    if (_T_1195) begin
      if (io_mem_s2_xcpt_ae_ld) begin
        if (r_req_dest) begin
          resp_valid_1 <= 1'h1;
        end else begin
          if (io_mem_resp_valid) begin
            if (_T_1200) begin
              resp_valid_1 <= r_req_dest;
            end else begin
              resp_valid_1 <= 1'h0;
            end
          end else begin
            resp_valid_1 <= 1'h0;
          end
        end
      end else begin
        if (io_mem_resp_valid) begin
          if (_T_1200) begin
            resp_valid_1 <= r_req_dest;
          end else begin
            resp_valid_1 <= 1'h0;
          end
        end else begin
          resp_valid_1 <= 1'h0;
        end
      end
    end else begin
      resp_valid_1 <= 1'h0;
    end
    if (_T_399) begin
      r_req_addr <= arb_io_out_bits_addr;
    end
    if (_T_399) begin
      r_req_dest <= arb_io_chosen;
    end
    if (_T_1195) begin
      if (io_mem_resp_valid) begin
        r_pte_ppn <= pte_ppn;
      end else begin
        if (_T_1186) begin
          if (pte_cache_hit) begin
            r_pte_ppn <= {{34'd0}, _T_521};
          end else begin
            if (_T_399) begin
              r_pte_ppn <= {{32'd0}, io_dpath_ptbr_ppn};
            end
          end
        end else begin
          if (_T_399) begin
            r_pte_ppn <= {{32'd0}, io_dpath_ptbr_ppn};
          end
        end
      end
    end else begin
      if (_T_1186) begin
        if (pte_cache_hit) begin
          r_pte_ppn <= {{34'd0}, _T_521};
        end else begin
          if (_T_399) begin
            r_pte_ppn <= {{32'd0}, io_dpath_ptbr_ppn};
          end
        end
      end else begin
        if (_T_399) begin
          r_pte_ppn <= {{32'd0}, io_dpath_ptbr_ppn};
        end
      end
    end
    if (_T_469) begin
      if (_T_491) begin
        _T_401 <= _T_494;
      end else begin
        _T_401 <= _T_497;
      end
    end
    if (reset) begin
      _T_404 <= 4'h0;
    end else begin
      if (_T_502) begin
        _T_404 <= 4'h0;
      end else begin
        if (_T_438) begin
          _T_404 <= _T_465;
        end
      end
    end
    if (_T_438) begin
      if (2'h0 == _T_462) begin
        _T_408_0 <= _GEN_0;
      end
    end
    if (_T_438) begin
      if (2'h1 == _T_462) begin
        _T_408_1 <= _GEN_0;
      end
    end
    if (_T_438) begin
      if (2'h2 == _T_462) begin
        _T_408_2 <= _GEN_0;
      end
    end
    if (_T_438) begin
      if (2'h3 == _T_462) begin
        _T_408_3 <= _GEN_0;
      end
    end
    if (_T_438) begin
      if (2'h0 == _T_462) begin
        _T_418_0 <= _GEN_1;
      end
    end
    if (_T_438) begin
      if (2'h1 == _T_462) begin
        _T_418_1 <= _GEN_1;
      end
    end
    if (_T_438) begin
      if (2'h2 == _T_462) begin
        _T_418_2 <= _GEN_1;
      end
    end
    if (_T_438) begin
      if (2'h3 == _T_462) begin
        _T_418_3 <= _GEN_1;
      end
    end
  end
endmodule
module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc
);
  wire [1:0] _T_4;
  wire  _T_6;
  wire [7:0] _T_7;
  wire  _T_9;
  wire [6:0] _T_12;
  wire [3:0] _T_13;
  wire [1:0] _T_14;
  wire  _T_15;
  wire  _T_16;
  wire [2:0] _T_18;
  wire [5:0] _T_19;
  wire [6:0] _T_20;
  wire [9:0] _T_21;
  wire [2:0] _T_25;
  wire [4:0] _T_26;
  wire [11:0] _T_27;
  wire [14:0] _T_28;
  wire [17:0] _T_29;
  wire [29:0] _T_30;
  wire [4:0] _T_38;
  wire [31:0] _T_40_bits;
  wire [1:0] _T_41;
  wire [2:0] _T_42;
  wire [4:0] _T_44;
  wire [7:0] _T_45;
  wire [2:0] _T_47;
  wire [4:0] _T_48;
  wire [11:0] _T_54;
  wire [12:0] _T_55;
  wire [15:0] _T_56;
  wire [27:0] _T_57;
  wire [31:0] _T_69_bits;
  wire [3:0] _T_75;
  wire [6:0] _T_76;
  wire [11:0] _T_85;
  wire [11:0] _T_86;
  wire [14:0] _T_87;
  wire [26:0] _T_88;
  wire [31:0] _T_100_bits;
  wire [26:0] _T_119;
  wire [31:0] _T_131_bits;
  wire [1:0] _T_139;
  wire [4:0] _T_154;
  wire [7:0] _T_156;
  wire [14:0] _T_157;
  wire [6:0] _T_158;
  wire [11:0] _T_159;
  wire [26:0] _T_160;
  wire [31:0] _T_172_bits;
  wire [2:0] _T_178;
  wire [4:0] _T_191;
  wire [7:0] _T_193;
  wire [14:0] _T_194;
  wire [7:0] _T_195;
  wire [12:0] _T_196;
  wire [27:0] _T_197;
  wire [31:0] _T_209_bits;
  wire [14:0] _T_235;
  wire [26:0] _T_238;
  wire [31:0] _T_250_bits;
  wire [14:0] _T_276;
  wire [26:0] _T_279;
  wire [31:0] _T_291_bits;
  wire  _T_292;
  wire [6:0] _T_296;
  wire [4:0] _T_297;
  wire [11:0] _T_298;
  wire [4:0] _T_299;
  wire [11:0] _T_303;
  wire [16:0] _T_304;
  wire [19:0] _T_305;
  wire [31:0] _T_306;
  wire [9:0] _T_319;
  wire  _T_320;
  wire [1:0] _T_321;
  wire  _T_323;
  wire  _T_324;
  wire  _T_325;
  wire [2:0] _T_326;
  wire [3:0] _T_328;
  wire [1:0] _T_329;
  wire [5:0] _T_330;
  wire [1:0] _T_331;
  wire [10:0] _T_332;
  wire [12:0] _T_333;
  wire [14:0] _T_334;
  wire [20:0] _T_335;
  wire  _T_336;
  wire [9:0] _T_358;
  wire  _T_380;
  wire [7:0] _T_402;
  wire [12:0] _T_405;
  wire [19:0] _T_406;
  wire [10:0] _T_407;
  wire [11:0] _T_408;
  wire [31:0] _T_409;
  wire [16:0] _T_430;
  wire [19:0] _T_431;
  wire [31:0] _T_432;
  wire  _T_449;
  wire [6:0] _T_452;
  wire [14:0] _T_457;
  wire [19:0] _T_460;
  wire [31:0] _T_461;
  wire [19:0] _T_462;
  wire [24:0] _T_464;
  wire [31:0] _T_465;
  wire  _T_476;
  wire  _T_479;
  wire  _T_480;
  wire [6:0] _T_492;
  wire [2:0] _T_497;
  wire [1:0] _T_498;
  wire [1:0] _T_503;
  wire [5:0] _T_504;
  wire [4:0] _T_505;
  wire [5:0] _T_506;
  wire [11:0] _T_507;
  wire [11:0] _T_511;
  wire [16:0] _T_512;
  wire [19:0] _T_513;
  wire [31:0] _T_514;
  wire [31:0] _T_523_bits;
  wire [4:0] _T_523_rd;
  wire [4:0] _T_523_rs2;
  wire [4:0] _T_523_rs3;
  wire [5:0] _T_526;
  wire [11:0] _T_535;
  wire [10:0] _T_536;
  wire [13:0] _T_537;
  wire [25:0] _T_538;
  wire [30:0] _GEN_0;
  wire [30:0] _T_555;
  wire [16:0] _T_572;
  wire [19:0] _T_573;
  wire [31:0] _T_574;
  wire [2:0] _T_585;
  wire  _T_587;
  wire [2:0] _T_588;
  wire  _T_590;
  wire [2:0] _T_591;
  wire  _T_593;
  wire [2:0] _T_594;
  wire  _T_596;
  wire [2:0] _T_597;
  wire  _T_599;
  wire [2:0] _T_600;
  wire  _T_602;
  wire [2:0] _T_603;
  wire  _T_605;
  wire [2:0] _T_606;
  wire  _T_609;
  wire [30:0] _T_612;
  wire [6:0] _T_616;
  wire [11:0] _T_626;
  wire [9:0] _T_627;
  wire [12:0] _T_628;
  wire [24:0] _T_629;
  wire [30:0] _GEN_1;
  wire [30:0] _T_630;
  wire [1:0] _T_631;
  wire  _T_633;
  wire [30:0] _T_634;
  wire  _T_636;
  wire [31:0] _T_637;
  wire  _T_639;
  wire [31:0] _T_640;
  wire [12:0] _T_743;
  wire [19:0] _T_744;
  wire [31:0] _T_747;
  wire [4:0] _T_762;
  wire [3:0] _T_768;
  wire [4:0] _T_769;
  wire [6:0] _T_770;
  wire [7:0] _T_771;
  wire [12:0] _T_772;
  wire  _T_773;
  wire [5:0] _T_789;
  wire [3:0] _T_810;
  wire  _T_826;
  wire [7:0] _T_828;
  wire [6:0] _T_829;
  wire [14:0] _T_830;
  wire [9:0] _T_831;
  wire [6:0] _T_832;
  wire [16:0] _T_833;
  wire [31:0] _T_834;
  wire [6:0] _T_916;
  wire [14:0] _T_917;
  wire [31:0] _T_921;
  wire [10:0] _T_938;
  wire [13:0] _T_939;
  wire [25:0] _T_940;
  wire [31:0] _T_946_bits;
  wire [4:0] _T_951;
  wire [3:0] _T_952;
  wire [8:0] _T_953;
  wire [11:0] _T_958;
  wire [13:0] _T_959;
  wire [16:0] _T_960;
  wire [28:0] _T_961;
  wire [31:0] _T_967_bits;
  wire [1:0] _T_968;
  wire [2:0] _T_970;
  wire [4:0] _T_972;
  wire [2:0] _T_973;
  wire [7:0] _T_974;
  wire [11:0] _T_979;
  wire [12:0] _T_980;
  wire [15:0] _T_981;
  wire [27:0] _T_982;
  wire [31:0] _T_988_bits;
  wire [27:0] _T_1003;
  wire [31:0] _T_1009_bits;
  wire [11:0] _T_1015;
  wire [9:0] _T_1016;
  wire [12:0] _T_1017;
  wire [24:0] _T_1018;
  wire [31:0] _T_1024_bits;
  wire [9:0] _T_1031;
  wire [12:0] _T_1032;
  wire [24:0] _T_1033;
  wire [31:0] _T_1039_bits;
  wire [24:0] _T_1048;
  wire [17:0] _T_1049;
  wire [24:0] _T_1051;
  wire  _T_1054;
  wire [24:0] _T_1055;
  wire [31:0] _T_1061_bits;
  wire  _T_1064;
  wire [31:0] _T_1065_bits;
  wire [4:0] _T_1065_rd;
  wire [4:0] _T_1065_rs1;
  wire [4:0] _T_1065_rs2;
  wire [4:0] _T_1065_rs3;
  wire [24:0] _T_1074;
  wire [24:0] _T_1077;
  wire [24:0] _T_1079;
  wire [24:0] _T_1083;
  wire [31:0] _T_1089_bits;
  wire [31:0] _T_1093_bits;
  wire [4:0] _T_1093_rd;
  wire [4:0] _T_1093_rs1;
  wire [31:0] _T_1095_bits;
  wire [4:0] _T_1095_rd;
  wire [4:0] _T_1095_rs1;
  wire [4:0] _T_1095_rs2;
  wire [4:0] _T_1095_rs3;
  wire [5:0] _T_1099;
  wire [8:0] _T_1100;
  wire [3:0] _T_1101;
  wire [4:0] _T_1110;
  wire [7:0] _T_1112;
  wire [14:0] _T_1113;
  wire [8:0] _T_1114;
  wire [13:0] _T_1115;
  wire [28:0] _T_1116;
  wire [31:0] _T_1122_bits;
  wire [1:0] _T_1123;
  wire [3:0] _T_1124;
  wire [5:0] _T_1126;
  wire [7:0] _T_1127;
  wire [2:0] _T_1128;
  wire [4:0] _T_1137;
  wire [7:0] _T_1139;
  wire [14:0] _T_1140;
  wire [7:0] _T_1141;
  wire [12:0] _T_1142;
  wire [27:0] _T_1143;
  wire [31:0] _T_1149_bits;
  wire [14:0] _T_1167;
  wire [27:0] _T_1170;
  wire [31:0] _T_1176_bits;
  wire [4:0] _T_1178;
  wire [4:0] _T_1179;
  wire [2:0] _T_1226;
  wire [4:0] _T_1227;
  wire  _T_1229;
  wire [31:0] _T_1230_bits;
  wire [4:0] _T_1230_rd;
  wire [4:0] _T_1230_rs1;
  wire [4:0] _T_1230_rs3;
  wire  _T_1232;
  wire [31:0] _T_1233_bits;
  wire [4:0] _T_1233_rd;
  wire [4:0] _T_1233_rs1;
  wire [4:0] _T_1233_rs3;
  wire  _T_1235;
  wire [31:0] _T_1236_bits;
  wire [4:0] _T_1236_rd;
  wire [4:0] _T_1236_rs1;
  wire [4:0] _T_1236_rs3;
  wire  _T_1238;
  wire [31:0] _T_1239_bits;
  wire [4:0] _T_1239_rd;
  wire [4:0] _T_1239_rs1;
  wire [4:0] _T_1239_rs3;
  wire  _T_1241;
  wire [31:0] _T_1242_bits;
  wire [4:0] _T_1242_rd;
  wire [4:0] _T_1242_rs1;
  wire [4:0] _T_1242_rs3;
  wire  _T_1244;
  wire [31:0] _T_1245_bits;
  wire [4:0] _T_1245_rd;
  wire [4:0] _T_1245_rs1;
  wire [4:0] _T_1245_rs3;
  wire  _T_1247;
  wire [31:0] _T_1248_bits;
  wire [4:0] _T_1248_rd;
  wire [4:0] _T_1248_rs1;
  wire [4:0] _T_1248_rs3;
  wire  _T_1250;
  wire [31:0] _T_1251_bits;
  wire [4:0] _T_1251_rd;
  wire [4:0] _T_1251_rs1;
  wire [4:0] _T_1251_rs2;
  wire [4:0] _T_1251_rs3;
  wire  _T_1253;
  wire [31:0] _T_1254_bits;
  wire [4:0] _T_1254_rd;
  wire [4:0] _T_1254_rs1;
  wire [4:0] _T_1254_rs2;
  wire [4:0] _T_1254_rs3;
  wire  _T_1256;
  wire [31:0] _T_1257_bits;
  wire [4:0] _T_1257_rd;
  wire [4:0] _T_1257_rs1;
  wire [4:0] _T_1257_rs2;
  wire [4:0] _T_1257_rs3;
  wire  _T_1259;
  wire [31:0] _T_1260_bits;
  wire [4:0] _T_1260_rd;
  wire [4:0] _T_1260_rs1;
  wire [4:0] _T_1260_rs2;
  wire [4:0] _T_1260_rs3;
  wire  _T_1262;
  wire [31:0] _T_1263_bits;
  wire [4:0] _T_1263_rd;
  wire [4:0] _T_1263_rs1;
  wire [4:0] _T_1263_rs2;
  wire [4:0] _T_1263_rs3;
  wire  _T_1265;
  wire [31:0] _T_1266_bits;
  wire [4:0] _T_1266_rd;
  wire [4:0] _T_1266_rs1;
  wire [4:0] _T_1266_rs2;
  wire [4:0] _T_1266_rs3;
  wire  _T_1268;
  wire [31:0] _T_1269_bits;
  wire [4:0] _T_1269_rd;
  wire [4:0] _T_1269_rs1;
  wire [4:0] _T_1269_rs2;
  wire [4:0] _T_1269_rs3;
  wire  _T_1271;
  wire [31:0] _T_1272_bits;
  wire [4:0] _T_1272_rd;
  wire [4:0] _T_1272_rs1;
  wire [4:0] _T_1272_rs2;
  wire [4:0] _T_1272_rs3;
  wire  _T_1274;
  wire [31:0] _T_1275_bits;
  wire [4:0] _T_1275_rd;
  wire [4:0] _T_1275_rs1;
  wire [4:0] _T_1275_rs2;
  wire [4:0] _T_1275_rs3;
  wire  _T_1277;
  wire [31:0] _T_1278_bits;
  wire [4:0] _T_1278_rd;
  wire [4:0] _T_1278_rs1;
  wire [4:0] _T_1278_rs2;
  wire [4:0] _T_1278_rs3;
  wire  _T_1280;
  wire [31:0] _T_1281_bits;
  wire [4:0] _T_1281_rd;
  wire [4:0] _T_1281_rs1;
  wire [4:0] _T_1281_rs2;
  wire [4:0] _T_1281_rs3;
  wire  _T_1283;
  wire [31:0] _T_1284_bits;
  wire [4:0] _T_1284_rd;
  wire [4:0] _T_1284_rs1;
  wire [4:0] _T_1284_rs2;
  wire [4:0] _T_1284_rs3;
  wire  _T_1286;
  wire [31:0] _T_1287_bits;
  wire [4:0] _T_1287_rd;
  wire [4:0] _T_1287_rs1;
  wire [4:0] _T_1287_rs2;
  wire [4:0] _T_1287_rs3;
  wire  _T_1289;
  wire [31:0] _T_1290_bits;
  wire [4:0] _T_1290_rd;
  wire [4:0] _T_1290_rs1;
  wire [4:0] _T_1290_rs2;
  wire [4:0] _T_1290_rs3;
  wire  _T_1292;
  wire [31:0] _T_1293_bits;
  wire [4:0] _T_1293_rd;
  wire [4:0] _T_1293_rs1;
  wire [4:0] _T_1293_rs2;
  wire [4:0] _T_1293_rs3;
  wire  _T_1295;
  wire [31:0] _T_1296_bits;
  wire [4:0] _T_1296_rd;
  wire [4:0] _T_1296_rs1;
  wire [4:0] _T_1296_rs2;
  wire [4:0] _T_1296_rs3;
  wire  _T_1298;
  wire [31:0] _T_1299_bits;
  wire [4:0] _T_1299_rd;
  wire [4:0] _T_1299_rs1;
  wire [4:0] _T_1299_rs2;
  wire [4:0] _T_1299_rs3;
  wire  _T_1301;
  wire [31:0] _T_1302_bits;
  wire [4:0] _T_1302_rd;
  wire [4:0] _T_1302_rs1;
  wire [4:0] _T_1302_rs2;
  wire [4:0] _T_1302_rs3;
  wire  _T_1304;
  wire [31:0] _T_1305_bits;
  wire [4:0] _T_1305_rd;
  wire [4:0] _T_1305_rs1;
  wire [4:0] _T_1305_rs2;
  wire [4:0] _T_1305_rs3;
  wire  _T_1307;
  wire [31:0] _T_1308_bits;
  wire [4:0] _T_1308_rd;
  wire [4:0] _T_1308_rs1;
  wire [4:0] _T_1308_rs2;
  wire [4:0] _T_1308_rs3;
  wire  _T_1310;
  wire [31:0] _T_1311_bits;
  wire [4:0] _T_1311_rd;
  wire [4:0] _T_1311_rs1;
  wire [4:0] _T_1311_rs2;
  wire [4:0] _T_1311_rs3;
  wire  _T_1313;
  wire [31:0] _T_1314_bits;
  wire [4:0] _T_1314_rd;
  wire [4:0] _T_1314_rs1;
  wire [4:0] _T_1314_rs2;
  wire [4:0] _T_1314_rs3;
  wire  _T_1316;
  wire [31:0] _T_1317_bits;
  wire [4:0] _T_1317_rd;
  wire [4:0] _T_1317_rs1;
  wire [4:0] _T_1317_rs2;
  wire [4:0] _T_1317_rs3;
  wire  _T_1319;
  wire [31:0] _T_1320_bits;
  wire [4:0] _T_1320_rd;
  wire [4:0] _T_1320_rs1;
  wire [4:0] _T_1320_rs2;
  wire [4:0] _T_1320_rs3;
  assign io_out_bits = _T_1320_bits;
  assign io_out_rd = _T_1320_rd;
  assign io_out_rs1 = _T_1320_rs1;
  assign io_out_rs2 = _T_1320_rs2;
  assign io_out_rs3 = _T_1320_rs3;
  assign io_rvc = _T_6;
  assign _T_4 = io_in[1:0];
  assign _T_6 = _T_4 != 2'h3;
  assign _T_7 = io_in[12:5];
  assign _T_9 = _T_7 != 8'h0;
  assign _T_12 = _T_9 ? 7'h13 : 7'h1f;
  assign _T_13 = io_in[10:7];
  assign _T_14 = io_in[12:11];
  assign _T_15 = io_in[5];
  assign _T_16 = io_in[6];
  assign _T_18 = {_T_16,2'h0};
  assign _T_19 = {_T_13,_T_14};
  assign _T_20 = {_T_19,_T_15};
  assign _T_21 = {_T_20,_T_18};
  assign _T_25 = io_in[4:2];
  assign _T_26 = {2'h1,_T_25};
  assign _T_27 = {_T_26,_T_12};
  assign _T_28 = {_T_21,5'h2};
  assign _T_29 = {_T_28,3'h0};
  assign _T_30 = {_T_29,_T_27};
  assign _T_38 = io_in[31:27];
  assign _T_40_bits = {{2'd0}, _T_30};
  assign _T_41 = io_in[6:5];
  assign _T_42 = io_in[12:10];
  assign _T_44 = {_T_41,_T_42};
  assign _T_45 = {_T_44,3'h0};
  assign _T_47 = io_in[9:7];
  assign _T_48 = {2'h1,_T_47};
  assign _T_54 = {_T_26,7'h7};
  assign _T_55 = {_T_45,_T_48};
  assign _T_56 = {_T_55,3'h3};
  assign _T_57 = {_T_56,_T_54};
  assign _T_69_bits = {{4'd0}, _T_57};
  assign _T_75 = {_T_15,_T_42};
  assign _T_76 = {_T_75,_T_18};
  assign _T_85 = {_T_26,7'h3};
  assign _T_86 = {_T_76,_T_48};
  assign _T_87 = {_T_86,3'h2};
  assign _T_88 = {_T_87,_T_85};
  assign _T_100_bits = {{5'd0}, _T_88};
  assign _T_119 = {_T_87,_T_54};
  assign _T_131_bits = {{5'd0}, _T_119};
  assign _T_139 = _T_76[6:5];
  assign _T_154 = _T_76[4:0];
  assign _T_156 = {3'h2,_T_154};
  assign _T_157 = {_T_156,7'h2f};
  assign _T_158 = {_T_139,_T_26};
  assign _T_159 = {_T_158,_T_48};
  assign _T_160 = {_T_159,_T_157};
  assign _T_172_bits = {{5'd0}, _T_160};
  assign _T_178 = _T_45[7:5];
  assign _T_191 = _T_45[4:0];
  assign _T_193 = {3'h3,_T_191};
  assign _T_194 = {_T_193,7'h27};
  assign _T_195 = {_T_178,_T_26};
  assign _T_196 = {_T_195,_T_48};
  assign _T_197 = {_T_196,_T_194};
  assign _T_209_bits = {{4'd0}, _T_197};
  assign _T_235 = {_T_156,7'h23};
  assign _T_238 = {_T_159,_T_235};
  assign _T_250_bits = {{5'd0}, _T_238};
  assign _T_276 = {_T_156,7'h27};
  assign _T_279 = {_T_159,_T_276};
  assign _T_291_bits = {{5'd0}, _T_279};
  assign _T_292 = io_in[12];
  assign _T_296 = _T_292 ? 7'h7f : 7'h0;
  assign _T_297 = io_in[6:2];
  assign _T_298 = {_T_296,_T_297};
  assign _T_299 = io_in[11:7];
  assign _T_303 = {_T_299,7'h13};
  assign _T_304 = {_T_298,_T_299};
  assign _T_305 = {_T_304,3'h0};
  assign _T_306 = {_T_305,_T_303};
  assign _T_319 = _T_292 ? 10'h3ff : 10'h0;
  assign _T_320 = io_in[8];
  assign _T_321 = io_in[10:9];
  assign _T_323 = io_in[7];
  assign _T_324 = io_in[2];
  assign _T_325 = io_in[11];
  assign _T_326 = io_in[5:3];
  assign _T_328 = {_T_326,1'h0};
  assign _T_329 = {_T_324,_T_325};
  assign _T_330 = {_T_329,_T_328};
  assign _T_331 = {_T_16,_T_323};
  assign _T_332 = {_T_319,_T_320};
  assign _T_333 = {_T_332,_T_321};
  assign _T_334 = {_T_333,_T_331};
  assign _T_335 = {_T_334,_T_330};
  assign _T_336 = _T_335[20];
  assign _T_358 = _T_335[10:1];
  assign _T_380 = _T_335[11];
  assign _T_402 = _T_335[19:12];
  assign _T_405 = {_T_402,5'h1};
  assign _T_406 = {_T_405,7'h6f};
  assign _T_407 = {_T_336,_T_358};
  assign _T_408 = {_T_407,_T_380};
  assign _T_409 = {_T_408,_T_406};
  assign _T_430 = {_T_298,5'h0};
  assign _T_431 = {_T_430,3'h0};
  assign _T_432 = {_T_431,_T_303};
  assign _T_449 = _T_298 != 12'h0;
  assign _T_452 = _T_449 ? 7'h37 : 7'h3f;
  assign _T_457 = _T_292 ? 15'h7fff : 15'h0;
  assign _T_460 = {_T_457,_T_297};
  assign _T_461 = {_T_460,12'h0};
  assign _T_462 = _T_461[31:12];
  assign _T_464 = {_T_462,_T_299};
  assign _T_465 = {_T_464,_T_452};
  assign _T_476 = _T_299 == 5'h0;
  assign _T_479 = _T_299 == 5'h2;
  assign _T_480 = _T_476 | _T_479;
  assign _T_492 = _T_449 ? 7'h13 : 7'h1f;
  assign _T_497 = _T_292 ? 3'h7 : 3'h0;
  assign _T_498 = io_in[4:3];
  assign _T_503 = {_T_324,_T_16};
  assign _T_504 = {_T_503,4'h0};
  assign _T_505 = {_T_497,_T_498};
  assign _T_506 = {_T_505,_T_15};
  assign _T_507 = {_T_506,_T_504};
  assign _T_511 = {_T_299,_T_492};
  assign _T_512 = {_T_507,_T_299};
  assign _T_513 = {_T_512,3'h0};
  assign _T_514 = {_T_513,_T_511};
  assign _T_523_bits = _T_480 ? _T_514 : _T_465;
  assign _T_523_rd = _T_480 ? _T_299 : _T_299;
  assign _T_523_rs2 = _T_480 ? _T_26 : _T_26;
  assign _T_523_rs3 = _T_480 ? _T_38 : _T_38;
  assign _T_526 = {_T_292,_T_297};
  assign _T_535 = {_T_48,7'h13};
  assign _T_536 = {_T_526,_T_48};
  assign _T_537 = {_T_536,3'h5};
  assign _T_538 = {_T_537,_T_535};
  assign _GEN_0 = {{5'd0}, _T_538};
  assign _T_555 = _GEN_0 | 31'h40000000;
  assign _T_572 = {_T_298,_T_48};
  assign _T_573 = {_T_572,3'h7};
  assign _T_574 = {_T_573,_T_535};
  assign _T_585 = {_T_292,_T_41};
  assign _T_587 = _T_585 == 3'h1;
  assign _T_588 = _T_587 ? 3'h4 : 3'h0;
  assign _T_590 = _T_585 == 3'h2;
  assign _T_591 = _T_590 ? 3'h6 : _T_588;
  assign _T_593 = _T_585 == 3'h3;
  assign _T_594 = _T_593 ? 3'h7 : _T_591;
  assign _T_596 = _T_585 == 3'h4;
  assign _T_597 = _T_596 ? 3'h0 : _T_594;
  assign _T_599 = _T_585 == 3'h5;
  assign _T_600 = _T_599 ? 3'h0 : _T_597;
  assign _T_602 = _T_585 == 3'h6;
  assign _T_603 = _T_602 ? 3'h2 : _T_600;
  assign _T_605 = _T_585 == 3'h7;
  assign _T_606 = _T_605 ? 3'h3 : _T_603;
  assign _T_609 = _T_41 == 2'h0;
  assign _T_612 = _T_609 ? 31'h40000000 : 31'h0;
  assign _T_616 = _T_292 ? 7'h3b : 7'h33;
  assign _T_626 = {_T_48,_T_616};
  assign _T_627 = {_T_26,_T_48};
  assign _T_628 = {_T_627,_T_606};
  assign _T_629 = {_T_628,_T_626};
  assign _GEN_1 = {{6'd0}, _T_629};
  assign _T_630 = _GEN_1 | _T_612;
  assign _T_631 = io_in[11:10];
  assign _T_633 = _T_631 == 2'h1;
  assign _T_634 = _T_633 ? _T_555 : {{5'd0}, _T_538};
  assign _T_636 = _T_631 == 2'h2;
  assign _T_637 = _T_636 ? _T_574 : {{1'd0}, _T_634};
  assign _T_639 = _T_631 == 2'h3;
  assign _T_640 = _T_639 ? {{1'd0}, _T_630} : _T_637;
  assign _T_743 = {_T_402,5'h0};
  assign _T_744 = {_T_743,7'h6f};
  assign _T_747 = {_T_408,_T_744};
  assign _T_762 = _T_292 ? 5'h1f : 5'h0;
  assign _T_768 = {_T_631,_T_498};
  assign _T_769 = {_T_768,1'h0};
  assign _T_770 = {_T_762,_T_41};
  assign _T_771 = {_T_770,_T_324};
  assign _T_772 = {_T_771,_T_769};
  assign _T_773 = _T_772[12];
  assign _T_789 = _T_772[10:5];
  assign _T_810 = _T_772[4:1];
  assign _T_826 = _T_772[11];
  assign _T_828 = {_T_826,7'h63};
  assign _T_829 = {3'h0,_T_810};
  assign _T_830 = {_T_829,_T_828};
  assign _T_831 = {5'h0,_T_48};
  assign _T_832 = {_T_773,_T_789};
  assign _T_833 = {_T_832,_T_831};
  assign _T_834 = {_T_833,_T_830};
  assign _T_916 = {3'h1,_T_810};
  assign _T_917 = {_T_916,_T_828};
  assign _T_921 = {_T_833,_T_917};
  assign _T_938 = {_T_526,_T_299};
  assign _T_939 = {_T_938,3'h1};
  assign _T_940 = {_T_939,_T_303};
  assign _T_946_bits = {{6'd0}, _T_940};
  assign _T_951 = {_T_41,3'h0};
  assign _T_952 = {_T_25,_T_292};
  assign _T_953 = {_T_952,_T_951};
  assign _T_958 = {_T_299,7'h7};
  assign _T_959 = {_T_953,5'h2};
  assign _T_960 = {_T_959,3'h3};
  assign _T_961 = {_T_960,_T_958};
  assign _T_967_bits = {{3'd0}, _T_961};
  assign _T_968 = io_in[3:2];
  assign _T_970 = io_in[6:4];
  assign _T_972 = {_T_970,2'h0};
  assign _T_973 = {_T_968,_T_292};
  assign _T_974 = {_T_973,_T_972};
  assign _T_979 = {_T_299,7'h3};
  assign _T_980 = {_T_974,5'h2};
  assign _T_981 = {_T_980,3'h2};
  assign _T_982 = {_T_981,_T_979};
  assign _T_988_bits = {{4'd0}, _T_982};
  assign _T_1003 = {_T_981,_T_958};
  assign _T_1009_bits = {{4'd0}, _T_1003};
  assign _T_1015 = {_T_299,7'h33};
  assign _T_1016 = {_T_297,5'h0};
  assign _T_1017 = {_T_1016,3'h0};
  assign _T_1018 = {_T_1017,_T_1015};
  assign _T_1024_bits = {{7'd0}, _T_1018};
  assign _T_1031 = {_T_297,_T_299};
  assign _T_1032 = {_T_1031,3'h0};
  assign _T_1033 = {_T_1032,_T_1015};
  assign _T_1039_bits = {{7'd0}, _T_1033};
  assign _T_1048 = {_T_1032,12'h67};
  assign _T_1049 = _T_1048[24:7];
  assign _T_1051 = {_T_1049,7'h1f};
  assign _T_1054 = _T_299 != 5'h0;
  assign _T_1055 = _T_1054 ? _T_1048 : _T_1051;
  assign _T_1061_bits = {{7'd0}, _T_1055};
  assign _T_1064 = _T_297 != 5'h0;
  assign _T_1065_bits = _T_1064 ? _T_1024_bits : _T_1061_bits;
  assign _T_1065_rd = _T_1064 ? _T_299 : 5'h0;
  assign _T_1065_rs1 = _T_1064 ? 5'h0 : _T_299;
  assign _T_1065_rs2 = _T_1064 ? _T_297 : _T_297;
  assign _T_1065_rs3 = _T_1064 ? _T_38 : _T_38;
  assign _T_1074 = {_T_1032,12'he7};
  assign _T_1077 = {_T_1049,7'h73};
  assign _T_1079 = _T_1077 | 25'h100000;
  assign _T_1083 = _T_1054 ? _T_1074 : _T_1079;
  assign _T_1089_bits = {{7'd0}, _T_1083};
  assign _T_1093_bits = _T_1064 ? _T_1039_bits : _T_1089_bits;
  assign _T_1093_rd = _T_1064 ? _T_299 : 5'h1;
  assign _T_1093_rs1 = _T_1064 ? _T_299 : _T_299;
  assign _T_1095_bits = _T_292 ? _T_1093_bits : _T_1065_bits;
  assign _T_1095_rd = _T_292 ? _T_1093_rd : _T_1065_rd;
  assign _T_1095_rs1 = _T_292 ? _T_1093_rs1 : _T_1065_rs1;
  assign _T_1095_rs2 = _T_292 ? _T_1065_rs2 : _T_1065_rs2;
  assign _T_1095_rs3 = _T_292 ? _T_1065_rs3 : _T_1065_rs3;
  assign _T_1099 = {_T_47,_T_42};
  assign _T_1100 = {_T_1099,3'h0};
  assign _T_1101 = _T_1100[8:5];
  assign _T_1110 = _T_1100[4:0];
  assign _T_1112 = {3'h3,_T_1110};
  assign _T_1113 = {_T_1112,7'h27};
  assign _T_1114 = {_T_1101,_T_297};
  assign _T_1115 = {_T_1114,5'h2};
  assign _T_1116 = {_T_1115,_T_1113};
  assign _T_1122_bits = {{3'd0}, _T_1116};
  assign _T_1123 = io_in[8:7];
  assign _T_1124 = io_in[12:9];
  assign _T_1126 = {_T_1123,_T_1124};
  assign _T_1127 = {_T_1126,2'h0};
  assign _T_1128 = _T_1127[7:5];
  assign _T_1137 = _T_1127[4:0];
  assign _T_1139 = {3'h2,_T_1137};
  assign _T_1140 = {_T_1139,7'h23};
  assign _T_1141 = {_T_1128,_T_297};
  assign _T_1142 = {_T_1141,5'h2};
  assign _T_1143 = {_T_1142,_T_1140};
  assign _T_1149_bits = {{4'd0}, _T_1143};
  assign _T_1167 = {_T_1139,7'h27};
  assign _T_1170 = {_T_1142,_T_1167};
  assign _T_1176_bits = {{4'd0}, _T_1170};
  assign _T_1178 = io_in[19:15];
  assign _T_1179 = io_in[24:20];
  assign _T_1226 = io_in[15:13];
  assign _T_1227 = {_T_4,_T_1226};
  assign _T_1229 = _T_1227 == 5'h1;
  assign _T_1230_bits = _T_1229 ? _T_69_bits : _T_40_bits;
  assign _T_1230_rd = _T_1229 ? _T_26 : _T_26;
  assign _T_1230_rs1 = _T_1229 ? _T_48 : 5'h2;
  assign _T_1230_rs3 = _T_1229 ? _T_38 : _T_38;
  assign _T_1232 = _T_1227 == 5'h2;
  assign _T_1233_bits = _T_1232 ? _T_100_bits : _T_1230_bits;
  assign _T_1233_rd = _T_1232 ? _T_26 : _T_1230_rd;
  assign _T_1233_rs1 = _T_1232 ? _T_48 : _T_1230_rs1;
  assign _T_1233_rs3 = _T_1232 ? _T_38 : _T_1230_rs3;
  assign _T_1235 = _T_1227 == 5'h3;
  assign _T_1236_bits = _T_1235 ? _T_131_bits : _T_1233_bits;
  assign _T_1236_rd = _T_1235 ? _T_26 : _T_1233_rd;
  assign _T_1236_rs1 = _T_1235 ? _T_48 : _T_1233_rs1;
  assign _T_1236_rs3 = _T_1235 ? _T_38 : _T_1233_rs3;
  assign _T_1238 = _T_1227 == 5'h4;
  assign _T_1239_bits = _T_1238 ? _T_172_bits : _T_1236_bits;
  assign _T_1239_rd = _T_1238 ? _T_26 : _T_1236_rd;
  assign _T_1239_rs1 = _T_1238 ? _T_48 : _T_1236_rs1;
  assign _T_1239_rs3 = _T_1238 ? _T_38 : _T_1236_rs3;
  assign _T_1241 = _T_1227 == 5'h5;
  assign _T_1242_bits = _T_1241 ? _T_209_bits : _T_1239_bits;
  assign _T_1242_rd = _T_1241 ? _T_26 : _T_1239_rd;
  assign _T_1242_rs1 = _T_1241 ? _T_48 : _T_1239_rs1;
  assign _T_1242_rs3 = _T_1241 ? _T_38 : _T_1239_rs3;
  assign _T_1244 = _T_1227 == 5'h6;
  assign _T_1245_bits = _T_1244 ? _T_250_bits : _T_1242_bits;
  assign _T_1245_rd = _T_1244 ? _T_26 : _T_1242_rd;
  assign _T_1245_rs1 = _T_1244 ? _T_48 : _T_1242_rs1;
  assign _T_1245_rs3 = _T_1244 ? _T_38 : _T_1242_rs3;
  assign _T_1247 = _T_1227 == 5'h7;
  assign _T_1248_bits = _T_1247 ? _T_291_bits : _T_1245_bits;
  assign _T_1248_rd = _T_1247 ? _T_26 : _T_1245_rd;
  assign _T_1248_rs1 = _T_1247 ? _T_48 : _T_1245_rs1;
  assign _T_1248_rs3 = _T_1247 ? _T_38 : _T_1245_rs3;
  assign _T_1250 = _T_1227 == 5'h8;
  assign _T_1251_bits = _T_1250 ? _T_306 : _T_1248_bits;
  assign _T_1251_rd = _T_1250 ? _T_299 : _T_1248_rd;
  assign _T_1251_rs1 = _T_1250 ? _T_299 : _T_1248_rs1;
  assign _T_1251_rs2 = _T_1250 ? _T_26 : _T_1248_rd;
  assign _T_1251_rs3 = _T_1250 ? _T_38 : _T_1248_rs3;
  assign _T_1253 = _T_1227 == 5'h9;
  assign _T_1254_bits = _T_1253 ? _T_409 : _T_1251_bits;
  assign _T_1254_rd = _T_1253 ? 5'h1 : _T_1251_rd;
  assign _T_1254_rs1 = _T_1253 ? _T_299 : _T_1251_rs1;
  assign _T_1254_rs2 = _T_1253 ? _T_26 : _T_1251_rs2;
  assign _T_1254_rs3 = _T_1253 ? _T_38 : _T_1251_rs3;
  assign _T_1256 = _T_1227 == 5'ha;
  assign _T_1257_bits = _T_1256 ? _T_432 : _T_1254_bits;
  assign _T_1257_rd = _T_1256 ? _T_299 : _T_1254_rd;
  assign _T_1257_rs1 = _T_1256 ? 5'h0 : _T_1254_rs1;
  assign _T_1257_rs2 = _T_1256 ? _T_26 : _T_1254_rs2;
  assign _T_1257_rs3 = _T_1256 ? _T_38 : _T_1254_rs3;
  assign _T_1259 = _T_1227 == 5'hb;
  assign _T_1260_bits = _T_1259 ? _T_523_bits : _T_1257_bits;
  assign _T_1260_rd = _T_1259 ? _T_523_rd : _T_1257_rd;
  assign _T_1260_rs1 = _T_1259 ? _T_523_rd : _T_1257_rs1;
  assign _T_1260_rs2 = _T_1259 ? _T_523_rs2 : _T_1257_rs2;
  assign _T_1260_rs3 = _T_1259 ? _T_523_rs3 : _T_1257_rs3;
  assign _T_1262 = _T_1227 == 5'hc;
  assign _T_1263_bits = _T_1262 ? _T_640 : _T_1260_bits;
  assign _T_1263_rd = _T_1262 ? _T_48 : _T_1260_rd;
  assign _T_1263_rs1 = _T_1262 ? _T_48 : _T_1260_rs1;
  assign _T_1263_rs2 = _T_1262 ? _T_26 : _T_1260_rs2;
  assign _T_1263_rs3 = _T_1262 ? _T_38 : _T_1260_rs3;
  assign _T_1265 = _T_1227 == 5'hd;
  assign _T_1266_bits = _T_1265 ? _T_747 : _T_1263_bits;
  assign _T_1266_rd = _T_1265 ? 5'h0 : _T_1263_rd;
  assign _T_1266_rs1 = _T_1265 ? _T_48 : _T_1263_rs1;
  assign _T_1266_rs2 = _T_1265 ? _T_26 : _T_1263_rs2;
  assign _T_1266_rs3 = _T_1265 ? _T_38 : _T_1263_rs3;
  assign _T_1268 = _T_1227 == 5'he;
  assign _T_1269_bits = _T_1268 ? _T_834 : _T_1266_bits;
  assign _T_1269_rd = _T_1268 ? _T_48 : _T_1266_rd;
  assign _T_1269_rs1 = _T_1268 ? _T_48 : _T_1266_rs1;
  assign _T_1269_rs2 = _T_1268 ? 5'h0 : _T_1266_rs2;
  assign _T_1269_rs3 = _T_1268 ? _T_38 : _T_1266_rs3;
  assign _T_1271 = _T_1227 == 5'hf;
  assign _T_1272_bits = _T_1271 ? _T_921 : _T_1269_bits;
  assign _T_1272_rd = _T_1271 ? 5'h0 : _T_1269_rd;
  assign _T_1272_rs1 = _T_1271 ? _T_48 : _T_1269_rs1;
  assign _T_1272_rs2 = _T_1271 ? 5'h0 : _T_1269_rs2;
  assign _T_1272_rs3 = _T_1271 ? _T_38 : _T_1269_rs3;
  assign _T_1274 = _T_1227 == 5'h10;
  assign _T_1275_bits = _T_1274 ? _T_946_bits : _T_1272_bits;
  assign _T_1275_rd = _T_1274 ? _T_299 : _T_1272_rd;
  assign _T_1275_rs1 = _T_1274 ? _T_299 : _T_1272_rs1;
  assign _T_1275_rs2 = _T_1274 ? _T_297 : _T_1272_rs2;
  assign _T_1275_rs3 = _T_1274 ? _T_38 : _T_1272_rs3;
  assign _T_1277 = _T_1227 == 5'h11;
  assign _T_1278_bits = _T_1277 ? _T_967_bits : _T_1275_bits;
  assign _T_1278_rd = _T_1277 ? _T_299 : _T_1275_rd;
  assign _T_1278_rs1 = _T_1277 ? 5'h2 : _T_1275_rs1;
  assign _T_1278_rs2 = _T_1277 ? _T_297 : _T_1275_rs2;
  assign _T_1278_rs3 = _T_1277 ? _T_38 : _T_1275_rs3;
  assign _T_1280 = _T_1227 == 5'h12;
  assign _T_1281_bits = _T_1280 ? _T_988_bits : _T_1278_bits;
  assign _T_1281_rd = _T_1280 ? _T_299 : _T_1278_rd;
  assign _T_1281_rs1 = _T_1280 ? 5'h2 : _T_1278_rs1;
  assign _T_1281_rs2 = _T_1280 ? _T_297 : _T_1278_rs2;
  assign _T_1281_rs3 = _T_1280 ? _T_38 : _T_1278_rs3;
  assign _T_1283 = _T_1227 == 5'h13;
  assign _T_1284_bits = _T_1283 ? _T_1009_bits : _T_1281_bits;
  assign _T_1284_rd = _T_1283 ? _T_299 : _T_1281_rd;
  assign _T_1284_rs1 = _T_1283 ? 5'h2 : _T_1281_rs1;
  assign _T_1284_rs2 = _T_1283 ? _T_297 : _T_1281_rs2;
  assign _T_1284_rs3 = _T_1283 ? _T_38 : _T_1281_rs3;
  assign _T_1286 = _T_1227 == 5'h14;
  assign _T_1287_bits = _T_1286 ? _T_1095_bits : _T_1284_bits;
  assign _T_1287_rd = _T_1286 ? _T_1095_rd : _T_1284_rd;
  assign _T_1287_rs1 = _T_1286 ? _T_1095_rs1 : _T_1284_rs1;
  assign _T_1287_rs2 = _T_1286 ? _T_1095_rs2 : _T_1284_rs2;
  assign _T_1287_rs3 = _T_1286 ? _T_1095_rs3 : _T_1284_rs3;
  assign _T_1289 = _T_1227 == 5'h15;
  assign _T_1290_bits = _T_1289 ? _T_1122_bits : _T_1287_bits;
  assign _T_1290_rd = _T_1289 ? _T_299 : _T_1287_rd;
  assign _T_1290_rs1 = _T_1289 ? 5'h2 : _T_1287_rs1;
  assign _T_1290_rs2 = _T_1289 ? _T_297 : _T_1287_rs2;
  assign _T_1290_rs3 = _T_1289 ? _T_38 : _T_1287_rs3;
  assign _T_1292 = _T_1227 == 5'h16;
  assign _T_1293_bits = _T_1292 ? _T_1149_bits : _T_1290_bits;
  assign _T_1293_rd = _T_1292 ? _T_299 : _T_1290_rd;
  assign _T_1293_rs1 = _T_1292 ? 5'h2 : _T_1290_rs1;
  assign _T_1293_rs2 = _T_1292 ? _T_297 : _T_1290_rs2;
  assign _T_1293_rs3 = _T_1292 ? _T_38 : _T_1290_rs3;
  assign _T_1295 = _T_1227 == 5'h17;
  assign _T_1296_bits = _T_1295 ? _T_1176_bits : _T_1293_bits;
  assign _T_1296_rd = _T_1295 ? _T_299 : _T_1293_rd;
  assign _T_1296_rs1 = _T_1295 ? 5'h2 : _T_1293_rs1;
  assign _T_1296_rs2 = _T_1295 ? _T_297 : _T_1293_rs2;
  assign _T_1296_rs3 = _T_1295 ? _T_38 : _T_1293_rs3;
  assign _T_1298 = _T_1227 == 5'h18;
  assign _T_1299_bits = _T_1298 ? io_in : _T_1296_bits;
  assign _T_1299_rd = _T_1298 ? _T_299 : _T_1296_rd;
  assign _T_1299_rs1 = _T_1298 ? _T_1178 : _T_1296_rs1;
  assign _T_1299_rs2 = _T_1298 ? _T_1179 : _T_1296_rs2;
  assign _T_1299_rs3 = _T_1298 ? _T_38 : _T_1296_rs3;
  assign _T_1301 = _T_1227 == 5'h19;
  assign _T_1302_bits = _T_1301 ? io_in : _T_1299_bits;
  assign _T_1302_rd = _T_1301 ? _T_299 : _T_1299_rd;
  assign _T_1302_rs1 = _T_1301 ? _T_1178 : _T_1299_rs1;
  assign _T_1302_rs2 = _T_1301 ? _T_1179 : _T_1299_rs2;
  assign _T_1302_rs3 = _T_1301 ? _T_38 : _T_1299_rs3;
  assign _T_1304 = _T_1227 == 5'h1a;
  assign _T_1305_bits = _T_1304 ? io_in : _T_1302_bits;
  assign _T_1305_rd = _T_1304 ? _T_299 : _T_1302_rd;
  assign _T_1305_rs1 = _T_1304 ? _T_1178 : _T_1302_rs1;
  assign _T_1305_rs2 = _T_1304 ? _T_1179 : _T_1302_rs2;
  assign _T_1305_rs3 = _T_1304 ? _T_38 : _T_1302_rs3;
  assign _T_1307 = _T_1227 == 5'h1b;
  assign _T_1308_bits = _T_1307 ? io_in : _T_1305_bits;
  assign _T_1308_rd = _T_1307 ? _T_299 : _T_1305_rd;
  assign _T_1308_rs1 = _T_1307 ? _T_1178 : _T_1305_rs1;
  assign _T_1308_rs2 = _T_1307 ? _T_1179 : _T_1305_rs2;
  assign _T_1308_rs3 = _T_1307 ? _T_38 : _T_1305_rs3;
  assign _T_1310 = _T_1227 == 5'h1c;
  assign _T_1311_bits = _T_1310 ? io_in : _T_1308_bits;
  assign _T_1311_rd = _T_1310 ? _T_299 : _T_1308_rd;
  assign _T_1311_rs1 = _T_1310 ? _T_1178 : _T_1308_rs1;
  assign _T_1311_rs2 = _T_1310 ? _T_1179 : _T_1308_rs2;
  assign _T_1311_rs3 = _T_1310 ? _T_38 : _T_1308_rs3;
  assign _T_1313 = _T_1227 == 5'h1d;
  assign _T_1314_bits = _T_1313 ? io_in : _T_1311_bits;
  assign _T_1314_rd = _T_1313 ? _T_299 : _T_1311_rd;
  assign _T_1314_rs1 = _T_1313 ? _T_1178 : _T_1311_rs1;
  assign _T_1314_rs2 = _T_1313 ? _T_1179 : _T_1311_rs2;
  assign _T_1314_rs3 = _T_1313 ? _T_38 : _T_1311_rs3;
  assign _T_1316 = _T_1227 == 5'h1e;
  assign _T_1317_bits = _T_1316 ? io_in : _T_1314_bits;
  assign _T_1317_rd = _T_1316 ? _T_299 : _T_1314_rd;
  assign _T_1317_rs1 = _T_1316 ? _T_1178 : _T_1314_rs1;
  assign _T_1317_rs2 = _T_1316 ? _T_1179 : _T_1314_rs2;
  assign _T_1317_rs3 = _T_1316 ? _T_38 : _T_1314_rs3;
  assign _T_1319 = _T_1227 == 5'h1f;
  assign _T_1320_bits = _T_1319 ? io_in : _T_1317_bits;
  assign _T_1320_rd = _T_1319 ? _T_299 : _T_1317_rd;
  assign _T_1320_rs1 = _T_1319 ? _T_1178 : _T_1317_rs1;
  assign _T_1320_rs2 = _T_1319 ? _T_1179 : _T_1317_rs2;
  assign _T_1320_rs3 = _T_1319 ? _T_38 : _T_1317_rs3;
endmodule
module IBuf(
  input         clock,
  input         reset,
  output        io_imem_ready,
  input         io_imem_valid,
  input         io_imem_bits_btb_valid,
  input         io_imem_bits_btb_bits_taken,
  input         io_imem_bits_btb_bits_bridx,
  input  [31:0] io_imem_bits_pc,
  input  [31:0] io_imem_bits_data,
  input         io_imem_bits_xcpt_pf_inst,
  input         io_imem_bits_xcpt_ae_inst,
  input         io_imem_bits_replay,
  input         io_kill,
  output [31:0] io_pc,
  input         io_inst_0_ready,
  output        io_inst_0_valid,
  output        io_inst_0_bits_xcpt0_pf_inst,
  output        io_inst_0_bits_xcpt0_ae_inst,
  output        io_inst_0_bits_xcpt1_pf_inst,
  output        io_inst_0_bits_xcpt1_ae_inst,
  output        io_inst_0_bits_replay,
  output        io_inst_0_bits_rvc,
  output [31:0] io_inst_0_bits_inst_bits,
  output [4:0]  io_inst_0_bits_inst_rd,
  output [4:0]  io_inst_0_bits_inst_rs1,
  output [4:0]  io_inst_0_bits_inst_rs2,
  output [4:0]  io_inst_0_bits_inst_rs3,
  output [31:0] io_inst_0_bits_raw
);
  reg  nBufValid;
  reg [31:0] _RAND_0;
  reg [31:0] buf_pc;
  reg [31:0] _RAND_1;
  reg [31:0] buf_data;
  reg [31:0] _RAND_2;
  reg  buf_xcpt_pf_inst;
  reg [31:0] _RAND_3;
  reg  buf_xcpt_ae_inst;
  reg [31:0] _RAND_4;
  reg  buf_replay;
  reg [31:0] _RAND_5;
  reg  ibufBTBHit;
  reg [31:0] _RAND_6;
  reg  ibufBTBResp_bridx;
  reg [31:0] _RAND_7;
  wire  pcWordBits;
  wire  _T_49;
  wire [1:0] _T_51;
  wire [1:0] _T_53;
  wire [1:0] _GEN_38;
  wire [2:0] _T_54;
  wire [2:0] _T_55;
  wire [1:0] nIC;
  wire [1:0] _GEN_39;
  wire [2:0] _T_56;
  wire [2:0] _T_57;
  wire [1:0] nICReady;
  wire [1:0] _T_59;
  wire [2:0] _T_60;
  wire [1:0] nValid;
  wire  _T_61;
  wire  _T_62;
  wire [2:0] _T_64;
  wire [2:0] _T_65;
  wire [1:0] _T_66;
  wire  _T_67;
  wire  _T_68;
  wire  _T_69;
  wire [2:0] _T_72;
  wire [2:0] _T_73;
  wire [1:0] _T_74;
  wire [1:0] _T_75;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  _T_85;
  wire [2:0] _T_86;
  wire [1:0] _T_87;
  wire [15:0] _T_91;
  wire [31:0] _T_92;
  wire [63:0] _T_93;
  wire [5:0] _GEN_46;
  wire [5:0] _T_94;
  wire [63:0] _T_95;
  wire [15:0] _T_96;
  wire [31:0] _T_98;
  wire [2:0] _GEN_47;
  wire [2:0] _T_99;
  wire [31:0] _GEN_48;
  wire [32:0] _T_100;
  wire [31:0] _T_101;
  wire [31:0] _T_102;
  wire [31:0] _T_103;
  wire [1:0] _GEN_49;
  wire [2:0] _T_104;
  wire [1:0] _T_105;
  wire [1:0] _GEN_3;
  wire [1:0] _GEN_9;
  wire [31:0] _GEN_20;
  wire [31:0] _GEN_21;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire [1:0] _GEN_30;
  wire [1:0] _GEN_36;
  wire [2:0] _T_108;
  wire [1:0] _T_109;
  wire [2:0] _T_110;
  wire [2:0] _T_111;
  wire [1:0] _T_112;
  wire [15:0] _T_113;
  wire [31:0] _T_114;
  wire [63:0] _T_115;
  wire [15:0] _T_116;
  wire [31:0] _T_117;
  wire [63:0] _T_118;
  wire [127:0] _T_119;
  wire [5:0] _GEN_52;
  wire [5:0] _T_120;
  wire [190:0] _GEN_53;
  wire [190:0] _T_121;
  wire [31:0] icData;
  wire [4:0] _GEN_54;
  wire [4:0] _T_124;
  wire [62:0] _T_125;
  wire [31:0] icMask;
  wire [31:0] _T_126;
  wire [31:0] _T_127;
  wire [31:0] _T_128;
  wire [31:0] inst;
  wire [3:0] _T_130;
  wire [4:0] _T_132;
  wire [4:0] _T_133;
  wire [3:0] _T_134;
  wire [1:0] valid;
  wire [1:0] _T_136;
  wire [2:0] _T_138;
  wire [2:0] _T_139;
  wire [1:0] bufMask;
  wire  _T_140;
  wire  xcpt_0_pf_inst;
  wire  xcpt_0_ae_inst;
  wire  _T_141;
  wire  xcpt_1_pf_inst;
  wire  xcpt_1_ae_inst;
  wire [1:0] _T_143;
  wire [1:0] _T_144;
  wire [1:0] _T_146;
  wire [1:0] _T_147;
  wire [1:0] ic_replay;
  wire [1:0] _T_149;
  wire [1:0] ibufBTBHitMask;
  wire  _T_152;
  wire  _T_154;
  wire  _T_155;
  wire  _T_156;
  wire  _T_157;
  wire  _T_158;
  wire  _T_160;
  wire [1:0] _T_161;
  wire [2:0] _T_162;
  wire [2:0] _T_163;
  wire [1:0] _T_164;
  wire [3:0] _T_166;
  wire [3:0] icBTBHitMask;
  wire [1:0] _T_168;
  wire [3:0] _GEN_56;
  wire [3:0] _T_170;
  wire [3:0] _GEN_57;
  wire [3:0] btbHitMask;
  wire  _T_176;
  wire [31:0] _T_177;
  wire [31:0] RVCExpander_io_in;
  wire [31:0] RVCExpander_io_out_bits;
  wire [4:0] RVCExpander_io_out_rd;
  wire [4:0] RVCExpander_io_out_rs1;
  wire [4:0] RVCExpander_io_out_rs2;
  wire [4:0] RVCExpander_io_out_rs3;
  wire  RVCExpander_io_rvc;
  wire [1:0] _T_179;
  wire  _T_180;
  wire  _T_182;
  wire [3:0] _T_183;
  wire  _T_184;
  wire [1:0] _T_186;
  wire  _T_187;
  wire [1:0] _T_188;
  wire  _T_189;
  wire  _T_190;
  wire  _T_191;
  wire  _T_192;
  wire [1:0] _T_193;
  wire  _T_194;
  wire [1:0] _T_198;
  wire  _T_199;
  wire  _T_200;
  wire  _T_206_pf_inst;
  wire  _T_206_ae_inst;
  wire [1:0] _T_207;
  wire  _T_209;
  wire  _T_210;
  wire  _T_211;
  wire  _T_212;
  wire [1:0] _T_224;
  wire  _T_230;
  wire  _T_231;
  wire  _T_243;
  wire [2:0] _T_248;
  wire [1:0] _T_249;
  wire [1:0] _T_250;
  wire [1:0] _GEN_37;
  RVCExpander RVCExpander (
    .io_in(RVCExpander_io_in),
    .io_out_bits(RVCExpander_io_out_bits),
    .io_out_rd(RVCExpander_io_out_rd),
    .io_out_rs1(RVCExpander_io_out_rs1),
    .io_out_rs2(RVCExpander_io_out_rs2),
    .io_out_rs3(RVCExpander_io_out_rs3),
    .io_rvc(RVCExpander_io_rvc)
  );
  assign io_imem_ready = _T_69;
  assign io_pc = _T_177;
  assign io_inst_0_valid = _T_212;
  assign io_inst_0_bits_xcpt0_pf_inst = xcpt_0_pf_inst;
  assign io_inst_0_bits_xcpt0_ae_inst = xcpt_0_ae_inst;
  assign io_inst_0_bits_xcpt1_pf_inst = _T_231;
  assign io_inst_0_bits_xcpt1_ae_inst = _T_230;
  assign io_inst_0_bits_replay = _T_192;
  assign io_inst_0_bits_rvc = RVCExpander_io_rvc;
  assign io_inst_0_bits_inst_bits = RVCExpander_io_out_bits;
  assign io_inst_0_bits_inst_rd = RVCExpander_io_out_rd;
  assign io_inst_0_bits_inst_rs1 = RVCExpander_io_out_rs1;
  assign io_inst_0_bits_inst_rs2 = RVCExpander_io_out_rs2;
  assign io_inst_0_bits_inst_rs3 = RVCExpander_io_out_rs3;
  assign io_inst_0_bits_raw = inst;
  assign pcWordBits = io_imem_bits_pc[1];
  assign _T_49 = io_imem_bits_btb_valid & io_imem_bits_btb_bits_taken;
  assign _T_51 = io_imem_bits_btb_bits_bridx + 1'h1;
  assign _T_53 = _T_49 ? _T_51 : 2'h2;
  assign _GEN_38 = {{1'd0}, pcWordBits};
  assign _T_54 = _T_53 - _GEN_38;
  assign _T_55 = $unsigned(_T_54);
  assign nIC = _T_55[1:0];
  assign _GEN_39 = {{1'd0}, nBufValid};
  assign _T_56 = _GEN_37 - _GEN_39;
  assign _T_57 = $unsigned(_T_56);
  assign nICReady = _T_57[1:0];
  assign _T_59 = io_imem_valid ? nIC : 2'h0;
  assign _T_60 = _T_59 + _GEN_39;
  assign nValid = _T_60[1:0];
  assign _T_61 = _GEN_37 >= _GEN_39;
  assign _T_62 = nICReady >= nIC;
  assign _T_64 = nIC - nICReady;
  assign _T_65 = $unsigned(_T_64);
  assign _T_66 = _T_65[1:0];
  assign _T_67 = 2'h1 >= _T_66;
  assign _T_68 = _T_62 | _T_67;
  assign _T_69 = _T_61 & _T_68;
  assign _T_72 = _GEN_39 - _GEN_37;
  assign _T_73 = $unsigned(_T_72);
  assign _T_74 = _T_73[1:0];
  assign _T_75 = _T_61 ? 2'h0 : _T_74;
  assign _T_77 = io_imem_valid & _T_61;
  assign _T_78 = nICReady < nIC;
  assign _T_79 = _T_77 & _T_78;
  assign _T_85 = _T_79 & _T_67;
  assign _T_86 = _GEN_38 + nICReady;
  assign _T_87 = _T_86[1:0];
  assign _T_91 = io_imem_bits_data[31:16];
  assign _T_92 = {_T_91,_T_91};
  assign _T_93 = {_T_92,io_imem_bits_data};
  assign _GEN_46 = {{4'd0}, _T_87};
  assign _T_94 = _GEN_46 << 4;
  assign _T_95 = _T_93 >> _T_94;
  assign _T_96 = _T_95[15:0];
  assign _T_98 = io_imem_bits_pc & 32'hfffffffc;
  assign _GEN_47 = {{1'd0}, nICReady};
  assign _T_99 = _GEN_47 << 1;
  assign _GEN_48 = {{29'd0}, _T_99};
  assign _T_100 = io_imem_bits_pc + _GEN_48;
  assign _T_101 = _T_100[31:0];
  assign _T_102 = _T_101 & 32'h3;
  assign _T_103 = _T_98 | _T_102;
  assign _GEN_49 = {{1'd0}, io_imem_bits_btb_bits_bridx};
  assign _T_104 = _GEN_49 + nICReady;
  assign _T_105 = _T_104[1:0];
  assign _GEN_3 = io_imem_bits_btb_valid ? _T_105 : {{1'd0}, ibufBTBResp_bridx};
  assign _GEN_9 = _T_85 ? _T_66 : _T_75;
  assign _GEN_20 = _T_85 ? _T_103 : buf_pc;
  assign _GEN_21 = _T_85 ? {{16'd0}, _T_96} : buf_data;
  assign _GEN_23 = _T_85 ? io_imem_bits_xcpt_pf_inst : buf_xcpt_pf_inst;
  assign _GEN_24 = _T_85 ? io_imem_bits_xcpt_ae_inst : buf_xcpt_ae_inst;
  assign _GEN_25 = _T_85 ? io_imem_bits_replay : buf_replay;
  assign _GEN_26 = _T_85 ? io_imem_bits_btb_valid : ibufBTBHit;
  assign _GEN_30 = _T_85 ? _GEN_3 : {{1'd0}, ibufBTBResp_bridx};
  assign _GEN_36 = io_kill ? 2'h0 : _GEN_9;
  assign _T_108 = 2'h2 + _GEN_39;
  assign _T_109 = _T_108[1:0];
  assign _T_110 = _T_109 - _GEN_38;
  assign _T_111 = $unsigned(_T_110);
  assign _T_112 = _T_111[1:0];
  assign _T_113 = io_imem_bits_data[15:0];
  assign _T_114 = {_T_113,_T_113};
  assign _T_115 = {io_imem_bits_data,_T_114};
  assign _T_116 = _T_115[63:48];
  assign _T_117 = {_T_116,_T_116};
  assign _T_118 = {_T_117,_T_117};
  assign _T_119 = {_T_118,_T_115};
  assign _GEN_52 = {{4'd0}, _T_112};
  assign _T_120 = _GEN_52 << 4;
  assign _GEN_53 = {{63'd0}, _T_119};
  assign _T_121 = _GEN_53 << _T_120;
  assign icData = _T_121[95:64];
  assign _GEN_54 = {{4'd0}, nBufValid};
  assign _T_124 = _GEN_54 << 4;
  assign _T_125 = 63'hffffffff << _T_124;
  assign icMask = _T_125[31:0];
  assign _T_126 = icData & icMask;
  assign _T_127 = ~ icMask;
  assign _T_128 = buf_data & _T_127;
  assign inst = _T_126 | _T_128;
  assign _T_130 = 4'h1 << nValid;
  assign _T_132 = _T_130 - 4'h1;
  assign _T_133 = $unsigned(_T_132);
  assign _T_134 = _T_133[3:0];
  assign valid = _T_134[1:0];
  assign _T_136 = 2'h1 << nBufValid;
  assign _T_138 = _T_136 - 2'h1;
  assign _T_139 = $unsigned(_T_138);
  assign bufMask = _T_139[1:0];
  assign _T_140 = bufMask[0];
  assign xcpt_0_pf_inst = _T_140 ? buf_xcpt_pf_inst : io_imem_bits_xcpt_pf_inst;
  assign xcpt_0_ae_inst = _T_140 ? buf_xcpt_ae_inst : io_imem_bits_xcpt_ae_inst;
  assign _T_141 = bufMask[1];
  assign xcpt_1_pf_inst = _T_141 ? buf_xcpt_pf_inst : io_imem_bits_xcpt_pf_inst;
  assign xcpt_1_ae_inst = _T_141 ? buf_xcpt_ae_inst : io_imem_bits_xcpt_ae_inst;
  assign _T_143 = buf_replay ? bufMask : 2'h0;
  assign _T_144 = ~ bufMask;
  assign _T_146 = io_imem_bits_replay ? _T_144 : 2'h0;
  assign _T_147 = _T_143 | _T_146;
  assign ic_replay = valid & _T_147;
  assign _T_149 = 2'h1 << ibufBTBResp_bridx;
  assign ibufBTBHitMask = ibufBTBHit ? _T_149 : 2'h0;
  assign _T_152 = io_imem_valid == 1'h0;
  assign _T_154 = io_imem_bits_btb_valid == 1'h0;
  assign _T_155 = _T_152 | _T_154;
  assign _T_156 = io_imem_bits_btb_bits_bridx >= pcWordBits;
  assign _T_157 = _T_155 | _T_156;
  assign _T_158 = _T_157 | reset;
  assign _T_160 = _T_158 == 1'h0;
  assign _T_161 = io_imem_bits_btb_bits_bridx + nBufValid;
  assign _T_162 = _T_161 - _GEN_38;
  assign _T_163 = $unsigned(_T_162);
  assign _T_164 = _T_163[1:0];
  assign _T_166 = 4'h1 << _T_164;
  assign icBTBHitMask = io_imem_bits_btb_valid ? _T_166 : 4'h0;
  assign _T_168 = ibufBTBHitMask & bufMask;
  assign _GEN_56 = {{2'd0}, _T_144};
  assign _T_170 = icBTBHitMask & _GEN_56;
  assign _GEN_57 = {{2'd0}, _T_168};
  assign btbHitMask = _GEN_57 | _T_170;
  assign _T_176 = nBufValid > 1'h0;
  assign _T_177 = _T_176 ? buf_pc : io_imem_bits_pc;
  assign RVCExpander_io_in = inst;
  assign _T_179 = ic_replay >> 1'h0;
  assign _T_180 = _T_179[0];
  assign _T_182 = RVCExpander_io_rvc == 1'h0;
  assign _T_183 = btbHitMask >> 1'h0;
  assign _T_184 = _T_183[0];
  assign _T_186 = 1'h0 + 1'h1;
  assign _T_187 = _T_186[0:0];
  assign _T_188 = ic_replay >> _T_187;
  assign _T_189 = _T_188[0];
  assign _T_190 = _T_184 | _T_189;
  assign _T_191 = _T_182 & _T_190;
  assign _T_192 = _T_180 | _T_191;
  assign _T_193 = valid >> 1'h0;
  assign _T_194 = _T_193[0];
  assign _T_198 = valid >> _T_187;
  assign _T_199 = _T_198[0];
  assign _T_200 = RVCExpander_io_rvc | _T_199;
  assign _T_206_pf_inst = _T_187 ? xcpt_1_pf_inst : xcpt_0_pf_inst;
  assign _T_206_ae_inst = _T_187 ? xcpt_1_ae_inst : xcpt_0_ae_inst;
  assign _T_207 = {_T_206_pf_inst,_T_206_ae_inst};
  assign _T_209 = _T_207 != 2'h0;
  assign _T_210 = _T_200 | _T_209;
  assign _T_211 = _T_210 | _T_192;
  assign _T_212 = _T_194 & _T_211;
  assign _T_224 = RVCExpander_io_rvc ? 2'h0 : _T_207;
  assign _T_230 = _T_224[0];
  assign _T_231 = _T_224[1];
  assign _T_243 = io_inst_0_ready & io_inst_0_valid;
  assign _T_248 = 2'h0 + 2'h2;
  assign _T_249 = _T_248[1:0];
  assign _T_250 = RVCExpander_io_rvc ? {{1'd0}, _T_187} : _T_249;
  assign _GEN_37 = _T_243 ? _T_250 : 2'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  nBufValid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  buf_pc = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  buf_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  buf_xcpt_pf_inst = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  buf_xcpt_ae_inst = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  buf_replay = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  ibufBTBHit = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  ibufBTBResp_bridx = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      nBufValid <= 1'h0;
    end else begin
      nBufValid <= _GEN_36[0];
    end
    if (_T_85) begin
      buf_pc <= _T_103;
    end
    if (_T_85) begin
      buf_data <= {{16'd0}, _T_96};
    end
    if (_T_85) begin
      buf_xcpt_pf_inst <= io_imem_bits_xcpt_pf_inst;
    end
    if (_T_85) begin
      buf_xcpt_ae_inst <= io_imem_bits_xcpt_ae_inst;
    end
    if (_T_85) begin
      buf_replay <= io_imem_bits_replay;
    end
    if (_T_85) begin
      ibufBTBHit <= io_imem_bits_btb_valid;
    end
    ibufBTBResp_bridx <= _GEN_30[0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_160) begin
          $fwrite(32'h80000002,"Assertion failed\n    at IBuf.scala:84 assert(!io.imem.valid || !io.imem.bits.btb.valid || io.imem.bits.btb.bits.bridx >= pcWordBits)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_160) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSRFile(
  input         clock,
  input         reset,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  input         io_hartid,
  input  [11:0] io_rw_addr,
  input  [2:0]  io_rw_cmd,
  output [31:0] io_rw_rdata,
  input  [31:0] io_rw_wdata,
  input  [11:0] io_decode_csr,
  output        io_decode_read_illegal,
  output        io_decode_write_illegal,
  output        io_decode_write_flush,
  output        io_decode_system_illegal,
  output        io_csr_stall,
  output        io_eret,
  output        io_singleStep,
  output        io_status_debug,
  output [31:0] io_status_isa,
  output [1:0]  io_status_dprv,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [26:0] io_status_zero2,
  output [1:0]  io_status_sxl,
  output [1:0]  io_status_uxl,
  output        io_status_sd_rv32,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_hpp,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [21:0] io_ptbr_ppn,
  output [31:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [31:0] io_cause,
  input  [31:0] io_pc,
  input  [31:0] io_badaddr,
  output [31:0] io_time,
  input         io_rocc_interrupt,
  output        io_interrupt,
  output [31:0] io_interrupt_cause,
  output        io_bp_0_control_action,
  output        io_bp_0_control_chain,
  output [1:0]  io_bp_0_control_tmatch,
  output        io_bp_0_control_m,
  output        io_bp_0_control_h,
  output        io_bp_0_control_s,
  output        io_bp_0_control_u,
  output        io_bp_0_control_x,
  output        io_bp_0_control_w,
  output        io_bp_0_control_r,
  output [31:0] io_bp_0_address,
  output        io_pmp_0_cfg_l,
  output [1:0]  io_pmp_0_cfg_a,
  output        io_pmp_0_cfg_x,
  output        io_pmp_0_cfg_w,
  output        io_pmp_0_cfg_r,
  output [29:0] io_pmp_0_addr,
  output [31:0] io_pmp_0_mask,
  output        io_pmp_1_cfg_l,
  output [1:0]  io_pmp_1_cfg_a,
  output        io_pmp_1_cfg_x,
  output        io_pmp_1_cfg_w,
  output        io_pmp_1_cfg_r,
  output [29:0] io_pmp_1_addr,
  output [31:0] io_pmp_1_mask,
  output        io_pmp_2_cfg_l,
  output [1:0]  io_pmp_2_cfg_a,
  output        io_pmp_2_cfg_x,
  output        io_pmp_2_cfg_w,
  output        io_pmp_2_cfg_r,
  output [29:0] io_pmp_2_addr,
  output [31:0] io_pmp_2_mask,
  output        io_pmp_3_cfg_l,
  output [1:0]  io_pmp_3_cfg_a,
  output        io_pmp_3_cfg_x,
  output        io_pmp_3_cfg_w,
  output        io_pmp_3_cfg_r,
  output [29:0] io_pmp_3_addr,
  output [31:0] io_pmp_3_mask,
  output        io_pmp_4_cfg_l,
  output [1:0]  io_pmp_4_cfg_a,
  output        io_pmp_4_cfg_x,
  output        io_pmp_4_cfg_w,
  output        io_pmp_4_cfg_r,
  output [29:0] io_pmp_4_addr,
  output [31:0] io_pmp_4_mask,
  output        io_pmp_5_cfg_l,
  output [1:0]  io_pmp_5_cfg_a,
  output        io_pmp_5_cfg_x,
  output        io_pmp_5_cfg_w,
  output        io_pmp_5_cfg_r,
  output [29:0] io_pmp_5_addr,
  output [31:0] io_pmp_5_mask,
  output        io_pmp_6_cfg_l,
  output [1:0]  io_pmp_6_cfg_a,
  output        io_pmp_6_cfg_x,
  output        io_pmp_6_cfg_w,
  output        io_pmp_6_cfg_r,
  output [29:0] io_pmp_6_addr,
  output [31:0] io_pmp_6_mask,
  output        io_pmp_7_cfg_l,
  output [1:0]  io_pmp_7_cfg_a,
  output        io_pmp_7_cfg_x,
  output        io_pmp_7_cfg_w,
  output        io_pmp_7_cfg_r,
  output [29:0] io_pmp_7_addr,
  output [31:0] io_pmp_7_mask
);
  reg [1:0] reg_mstatus_prv;
  reg [31:0] _RAND_0;
  reg [26:0] reg_mstatus_zero2;
  reg [31:0] _RAND_1;
  reg [7:0] reg_mstatus_zero1;
  reg [31:0] _RAND_2;
  reg  reg_mstatus_tsr;
  reg [31:0] _RAND_3;
  reg  reg_mstatus_tw;
  reg [31:0] _RAND_4;
  reg  reg_mstatus_tvm;
  reg [31:0] _RAND_5;
  reg  reg_mstatus_mxr;
  reg [31:0] _RAND_6;
  reg  reg_mstatus_sum;
  reg [31:0] _RAND_7;
  reg  reg_mstatus_mprv;
  reg [31:0] _RAND_8;
  reg [1:0] reg_mstatus_xs;
  reg [31:0] _RAND_9;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] _RAND_10;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] _RAND_11;
  reg [1:0] reg_mstatus_hpp;
  reg [31:0] _RAND_12;
  reg  reg_mstatus_spp;
  reg [31:0] _RAND_13;
  reg  reg_mstatus_mpie;
  reg [31:0] _RAND_14;
  reg  reg_mstatus_hpie;
  reg [31:0] _RAND_15;
  reg  reg_mstatus_spie;
  reg [31:0] _RAND_16;
  reg  reg_mstatus_upie;
  reg [31:0] _RAND_17;
  reg  reg_mstatus_mie;
  reg [31:0] _RAND_18;
  reg  reg_mstatus_hie;
  reg [31:0] _RAND_19;
  reg  reg_mstatus_sie;
  reg [31:0] _RAND_20;
  reg  reg_mstatus_uie;
  reg [31:0] _RAND_21;
  reg [1:0] reg_dcsr_xdebugver;
  reg [31:0] _RAND_22;
  reg [1:0] reg_dcsr_zero4;
  reg [31:0] _RAND_23;
  reg [11:0] reg_dcsr_zero3;
  reg [31:0] _RAND_24;
  reg  reg_dcsr_ebreakm;
  reg [31:0] _RAND_25;
  reg  reg_dcsr_ebreakh;
  reg [31:0] _RAND_26;
  reg  reg_dcsr_ebreaks;
  reg [31:0] _RAND_27;
  reg  reg_dcsr_ebreaku;
  reg [31:0] _RAND_28;
  reg  reg_dcsr_zero2;
  reg [31:0] _RAND_29;
  reg  reg_dcsr_stopcycle;
  reg [31:0] _RAND_30;
  reg  reg_dcsr_stoptime;
  reg [31:0] _RAND_31;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] _RAND_32;
  reg [2:0] reg_dcsr_zero1;
  reg [31:0] _RAND_33;
  reg  reg_dcsr_step;
  reg [31:0] _RAND_34;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] _RAND_35;
  reg  reg_debugint;
  reg [31:0] _RAND_36;
  reg  reg_debug;
  reg [31:0] _RAND_37;
  reg [31:0] reg_dpc;
  reg [31:0] _RAND_38;
  reg [31:0] reg_dscratch;
  reg [31:0] _RAND_39;
  reg  reg_singleStepped;
  reg [31:0] _RAND_40;
  reg  reg_tselect;
  reg [31:0] _RAND_41;
  reg [3:0] reg_bp_0_control_ttype;
  reg [31:0] _RAND_42;
  reg  reg_bp_0_control_dmode;
  reg [31:0] _RAND_43;
  reg [5:0] reg_bp_0_control_maskmax;
  reg [31:0] _RAND_44;
  reg [7:0] reg_bp_0_control_reserved;
  reg [31:0] _RAND_45;
  reg  reg_bp_0_control_action;
  reg [31:0] _RAND_46;
  reg  reg_bp_0_control_chain;
  reg [31:0] _RAND_47;
  reg [1:0] reg_bp_0_control_zero;
  reg [31:0] _RAND_48;
  reg [1:0] reg_bp_0_control_tmatch;
  reg [31:0] _RAND_49;
  reg  reg_bp_0_control_m;
  reg [31:0] _RAND_50;
  reg  reg_bp_0_control_h;
  reg [31:0] _RAND_51;
  reg  reg_bp_0_control_s;
  reg [31:0] _RAND_52;
  reg  reg_bp_0_control_u;
  reg [31:0] _RAND_53;
  reg  reg_bp_0_control_x;
  reg [31:0] _RAND_54;
  reg  reg_bp_0_control_w;
  reg [31:0] _RAND_55;
  reg  reg_bp_0_control_r;
  reg [31:0] _RAND_56;
  reg [31:0] reg_bp_0_address;
  reg [31:0] _RAND_57;
  reg [3:0] reg_bp_1_control_ttype;
  reg [31:0] _RAND_58;
  reg  reg_bp_1_control_dmode;
  reg [31:0] _RAND_59;
  reg [5:0] reg_bp_1_control_maskmax;
  reg [31:0] _RAND_60;
  reg [7:0] reg_bp_1_control_reserved;
  reg [31:0] _RAND_61;
  reg  reg_bp_1_control_action;
  reg [31:0] _RAND_62;
  reg  reg_bp_1_control_chain;
  reg [31:0] _RAND_63;
  reg [1:0] reg_bp_1_control_zero;
  reg [31:0] _RAND_64;
  reg [1:0] reg_bp_1_control_tmatch;
  reg [31:0] _RAND_65;
  reg  reg_bp_1_control_m;
  reg [31:0] _RAND_66;
  reg  reg_bp_1_control_h;
  reg [31:0] _RAND_67;
  reg  reg_bp_1_control_s;
  reg [31:0] _RAND_68;
  reg  reg_bp_1_control_u;
  reg [31:0] _RAND_69;
  reg  reg_bp_1_control_x;
  reg [31:0] _RAND_70;
  reg  reg_bp_1_control_w;
  reg [31:0] _RAND_71;
  reg  reg_bp_1_control_r;
  reg [31:0] _RAND_72;
  reg [31:0] reg_bp_1_address;
  reg [31:0] _RAND_73;
  reg  reg_pmp_0_cfg_l;
  reg [31:0] _RAND_74;
  reg [1:0] reg_pmp_0_cfg_res;
  reg [31:0] _RAND_75;
  reg [1:0] reg_pmp_0_cfg_a;
  reg [31:0] _RAND_76;
  reg  reg_pmp_0_cfg_x;
  reg [31:0] _RAND_77;
  reg  reg_pmp_0_cfg_w;
  reg [31:0] _RAND_78;
  reg  reg_pmp_0_cfg_r;
  reg [31:0] _RAND_79;
  reg [29:0] reg_pmp_0_addr;
  reg [31:0] _RAND_80;
  reg  reg_pmp_1_cfg_l;
  reg [31:0] _RAND_81;
  reg [1:0] reg_pmp_1_cfg_res;
  reg [31:0] _RAND_82;
  reg [1:0] reg_pmp_1_cfg_a;
  reg [31:0] _RAND_83;
  reg  reg_pmp_1_cfg_x;
  reg [31:0] _RAND_84;
  reg  reg_pmp_1_cfg_w;
  reg [31:0] _RAND_85;
  reg  reg_pmp_1_cfg_r;
  reg [31:0] _RAND_86;
  reg [29:0] reg_pmp_1_addr;
  reg [31:0] _RAND_87;
  reg  reg_pmp_2_cfg_l;
  reg [31:0] _RAND_88;
  reg [1:0] reg_pmp_2_cfg_res;
  reg [31:0] _RAND_89;
  reg [1:0] reg_pmp_2_cfg_a;
  reg [31:0] _RAND_90;
  reg  reg_pmp_2_cfg_x;
  reg [31:0] _RAND_91;
  reg  reg_pmp_2_cfg_w;
  reg [31:0] _RAND_92;
  reg  reg_pmp_2_cfg_r;
  reg [31:0] _RAND_93;
  reg [29:0] reg_pmp_2_addr;
  reg [31:0] _RAND_94;
  reg  reg_pmp_3_cfg_l;
  reg [31:0] _RAND_95;
  reg [1:0] reg_pmp_3_cfg_res;
  reg [31:0] _RAND_96;
  reg [1:0] reg_pmp_3_cfg_a;
  reg [31:0] _RAND_97;
  reg  reg_pmp_3_cfg_x;
  reg [31:0] _RAND_98;
  reg  reg_pmp_3_cfg_w;
  reg [31:0] _RAND_99;
  reg  reg_pmp_3_cfg_r;
  reg [31:0] _RAND_100;
  reg [29:0] reg_pmp_3_addr;
  reg [31:0] _RAND_101;
  reg  reg_pmp_4_cfg_l;
  reg [31:0] _RAND_102;
  reg [1:0] reg_pmp_4_cfg_res;
  reg [31:0] _RAND_103;
  reg [1:0] reg_pmp_4_cfg_a;
  reg [31:0] _RAND_104;
  reg  reg_pmp_4_cfg_x;
  reg [31:0] _RAND_105;
  reg  reg_pmp_4_cfg_w;
  reg [31:0] _RAND_106;
  reg  reg_pmp_4_cfg_r;
  reg [31:0] _RAND_107;
  reg [29:0] reg_pmp_4_addr;
  reg [31:0] _RAND_108;
  reg  reg_pmp_5_cfg_l;
  reg [31:0] _RAND_109;
  reg [1:0] reg_pmp_5_cfg_res;
  reg [31:0] _RAND_110;
  reg [1:0] reg_pmp_5_cfg_a;
  reg [31:0] _RAND_111;
  reg  reg_pmp_5_cfg_x;
  reg [31:0] _RAND_112;
  reg  reg_pmp_5_cfg_w;
  reg [31:0] _RAND_113;
  reg  reg_pmp_5_cfg_r;
  reg [31:0] _RAND_114;
  reg [29:0] reg_pmp_5_addr;
  reg [31:0] _RAND_115;
  reg  reg_pmp_6_cfg_l;
  reg [31:0] _RAND_116;
  reg [1:0] reg_pmp_6_cfg_res;
  reg [31:0] _RAND_117;
  reg [1:0] reg_pmp_6_cfg_a;
  reg [31:0] _RAND_118;
  reg  reg_pmp_6_cfg_x;
  reg [31:0] _RAND_119;
  reg  reg_pmp_6_cfg_w;
  reg [31:0] _RAND_120;
  reg  reg_pmp_6_cfg_r;
  reg [31:0] _RAND_121;
  reg [29:0] reg_pmp_6_addr;
  reg [31:0] _RAND_122;
  reg  reg_pmp_7_cfg_l;
  reg [31:0] _RAND_123;
  reg [1:0] reg_pmp_7_cfg_res;
  reg [31:0] _RAND_124;
  reg [1:0] reg_pmp_7_cfg_a;
  reg [31:0] _RAND_125;
  reg  reg_pmp_7_cfg_x;
  reg [31:0] _RAND_126;
  reg  reg_pmp_7_cfg_w;
  reg [31:0] _RAND_127;
  reg  reg_pmp_7_cfg_r;
  reg [31:0] _RAND_128;
  reg [29:0] reg_pmp_7_addr;
  reg [31:0] _RAND_129;
  reg [31:0] reg_mie;
  reg [31:0] _RAND_130;
  reg [31:0] reg_mideleg;
  reg [31:0] _RAND_131;
  reg  reg_mip_zero2;
  reg [31:0] _RAND_132;
  reg  reg_mip_debug;
  reg [31:0] _RAND_133;
  reg  reg_mip_zero1;
  reg [31:0] _RAND_134;
  reg  reg_mip_meip;
  reg [31:0] _RAND_135;
  reg  reg_mip_heip;
  reg [31:0] _RAND_136;
  reg  reg_mip_seip;
  reg [31:0] _RAND_137;
  reg  reg_mip_ueip;
  reg [31:0] _RAND_138;
  reg  reg_mip_mtip;
  reg [31:0] _RAND_139;
  reg  reg_mip_htip;
  reg [31:0] _RAND_140;
  reg  reg_mip_stip;
  reg [31:0] _RAND_141;
  reg  reg_mip_utip;
  reg [31:0] _RAND_142;
  reg  reg_mip_msip;
  reg [31:0] _RAND_143;
  reg  reg_mip_hsip;
  reg [31:0] _RAND_144;
  reg  reg_mip_ssip;
  reg [31:0] _RAND_145;
  reg  reg_mip_usip;
  reg [31:0] _RAND_146;
  reg [31:0] reg_mepc;
  reg [31:0] _RAND_147;
  reg [31:0] reg_mcause;
  reg [31:0] _RAND_148;
  reg [31:0] reg_mbadaddr;
  reg [31:0] _RAND_149;
  reg [31:0] reg_mscratch;
  reg [31:0] _RAND_150;
  reg [31:0] reg_mtvec;
  reg [31:0] _RAND_151;
  reg [31:0] reg_mcounteren;
  reg [31:0] _RAND_152;
  reg [21:0] reg_sptbr_ppn;
  reg [31:0] _RAND_153;
  reg  reg_wfi;
  reg [31:0] _RAND_154;
  reg [5:0] _T_248;
  reg [31:0] _RAND_155;
  wire [5:0] _GEN_0;
  wire [6:0] _T_249;
  reg [57:0] _T_252;
  reg [63:0] _RAND_156;
  wire  _T_253;
  wire [58:0] _T_255;
  wire [57:0] _T_256;
  wire [57:0] _GEN_35;
  wire [63:0] _T_257;
  reg [5:0] _T_261;
  reg [31:0] _RAND_157;
  wire [6:0] _T_262;
  reg [57:0] _T_265;
  reg [63:0] _RAND_158;
  wire  _T_266;
  wire [58:0] _T_268;
  wire [57:0] _T_269;
  wire [57:0] _GEN_36;
  wire [63:0] _T_270;
  wire  _T_273;
  wire [31:0] hpm_mask;
  wire [1:0] _T_282;
  wire [1:0] _T_283;
  wire [3:0] _T_284;
  wire [1:0] _T_285;
  wire [1:0] _T_286;
  wire [3:0] _T_287;
  wire [7:0] _T_288;
  wire [1:0] _T_289;
  wire [1:0] _T_290;
  wire [3:0] _T_291;
  wire [1:0] _T_292;
  wire [1:0] _T_293;
  wire [3:0] _T_294;
  wire [7:0] _T_295;
  wire [15:0] _T_296;
  wire [15:0] read_mip;
  wire [31:0] _GEN_1;
  wire [31:0] pending_interrupts;
  wire [14:0] _GEN_2;
  wire [14:0] d_interrupts;
  wire  _T_298;
  wire  _T_300;
  wire  _T_301;
  wire  _T_302;
  wire [31:0] _T_303;
  wire [31:0] _T_304;
  wire [31:0] m_interrupts;
  wire  _T_307;
  wire  _T_309;
  wire  _T_312;
  wire  _T_313;
  wire  _T_314;
  wire [31:0] _T_315;
  wire [31:0] s_interrupts;
  wire [31:0] _T_319;
  wire [31:0] _T_320;
  wire [63:0] _T_321;
  wire [31:0] _T_323;
  wire [31:0] _T_324;
  wire [63:0] _T_325;
  wire [31:0] _T_327;
  wire [31:0] _T_329;
  wire [31:0] _T_332;
  wire [63:0] _T_333;
  wire  _T_335;
  wire  _T_337;
  wire  _T_339;
  wire  _T_340;
  wire  anyInterrupt;
  wire [127:0] _T_341;
  wire [191:0] _T_342;
  wire [63:0] _T_343;
  wire [127:0] _T_344;
  wire  _T_346;
  wire [31:0] _T_347;
  wire [31:0] _T_348;
  wire  _T_350;
  wire [15:0] _T_351;
  wire [15:0] _T_352;
  wire  _T_354;
  wire [7:0] _T_355;
  wire [7:0] _T_356;
  wire  _T_358;
  wire [3:0] _T_359;
  wire [3:0] _T_360;
  wire  _T_362;
  wire  _T_363;
  wire  _T_365;
  wire  _T_367;
  wire [1:0] _T_368;
  wire [1:0] _T_369;
  wire  _T_370;
  wire  _T_372;
  wire  _T_374;
  wire [1:0] _T_375;
  wire [1:0] _T_376;
  wire [1:0] _T_377;
  wire [2:0] _T_378;
  wire [3:0] _T_379;
  wire [3:0] _T_380;
  wire  _T_382;
  wire  _T_383;
  wire  _T_385;
  wire  _T_387;
  wire [1:0] _T_388;
  wire [1:0] _T_389;
  wire  _T_390;
  wire  _T_392;
  wire  _T_394;
  wire [1:0] _T_395;
  wire [1:0] _T_396;
  wire [1:0] _T_397;
  wire [2:0] _T_398;
  wire [2:0] _T_399;
  wire [3:0] _T_400;
  wire [7:0] _T_401;
  wire [7:0] _T_402;
  wire  _T_404;
  wire [3:0] _T_405;
  wire [3:0] _T_406;
  wire  _T_408;
  wire  _T_409;
  wire  _T_411;
  wire  _T_413;
  wire [1:0] _T_414;
  wire [1:0] _T_415;
  wire  _T_416;
  wire  _T_418;
  wire  _T_420;
  wire [1:0] _T_421;
  wire [1:0] _T_422;
  wire [1:0] _T_423;
  wire [2:0] _T_424;
  wire [3:0] _T_425;
  wire [3:0] _T_426;
  wire  _T_428;
  wire  _T_429;
  wire  _T_431;
  wire  _T_433;
  wire [1:0] _T_434;
  wire [1:0] _T_435;
  wire  _T_436;
  wire  _T_438;
  wire  _T_440;
  wire [1:0] _T_441;
  wire [1:0] _T_442;
  wire [1:0] _T_443;
  wire [2:0] _T_444;
  wire [2:0] _T_445;
  wire [3:0] _T_446;
  wire [3:0] _T_447;
  wire [4:0] _T_448;
  wire [15:0] _T_449;
  wire [15:0] _T_450;
  wire  _T_452;
  wire [7:0] _T_453;
  wire [7:0] _T_454;
  wire  _T_456;
  wire [3:0] _T_457;
  wire [3:0] _T_458;
  wire  _T_460;
  wire  _T_461;
  wire  _T_463;
  wire  _T_465;
  wire [1:0] _T_466;
  wire [1:0] _T_467;
  wire  _T_468;
  wire  _T_470;
  wire  _T_472;
  wire [1:0] _T_473;
  wire [1:0] _T_474;
  wire [1:0] _T_475;
  wire [2:0] _T_476;
  wire [3:0] _T_477;
  wire [3:0] _T_478;
  wire  _T_480;
  wire  _T_481;
  wire  _T_483;
  wire  _T_485;
  wire [1:0] _T_486;
  wire [1:0] _T_487;
  wire  _T_488;
  wire  _T_490;
  wire  _T_492;
  wire [1:0] _T_493;
  wire [1:0] _T_494;
  wire [1:0] _T_495;
  wire [2:0] _T_496;
  wire [2:0] _T_497;
  wire [3:0] _T_498;
  wire [7:0] _T_499;
  wire [7:0] _T_500;
  wire  _T_502;
  wire [3:0] _T_503;
  wire [3:0] _T_504;
  wire  _T_506;
  wire  _T_507;
  wire  _T_509;
  wire  _T_511;
  wire [1:0] _T_512;
  wire [1:0] _T_513;
  wire  _T_514;
  wire  _T_516;
  wire  _T_518;
  wire [1:0] _T_519;
  wire [1:0] _T_520;
  wire [1:0] _T_521;
  wire [2:0] _T_522;
  wire [3:0] _T_523;
  wire [3:0] _T_524;
  wire  _T_526;
  wire  _T_527;
  wire  _T_529;
  wire  _T_531;
  wire [1:0] _T_532;
  wire [1:0] _T_533;
  wire  _T_534;
  wire  _T_536;
  wire  _T_538;
  wire [1:0] _T_539;
  wire [1:0] _T_540;
  wire [1:0] _T_541;
  wire [2:0] _T_542;
  wire [2:0] _T_543;
  wire [3:0] _T_544;
  wire [3:0] _T_545;
  wire [4:0] _T_546;
  wire [4:0] _T_547;
  wire [5:0] _T_548;
  wire [63:0] _T_549;
  wire [63:0] _T_550;
  wire  _T_552;
  wire [31:0] _T_553;
  wire [31:0] _T_554;
  wire  _T_556;
  wire [15:0] _T_557;
  wire [15:0] _T_558;
  wire  _T_560;
  wire [7:0] _T_561;
  wire [7:0] _T_562;
  wire  _T_564;
  wire [3:0] _T_565;
  wire [3:0] _T_566;
  wire  _T_568;
  wire  _T_569;
  wire  _T_571;
  wire  _T_573;
  wire [1:0] _T_574;
  wire [1:0] _T_575;
  wire  _T_576;
  wire  _T_578;
  wire  _T_580;
  wire [1:0] _T_581;
  wire [1:0] _T_582;
  wire [1:0] _T_583;
  wire [2:0] _T_584;
  wire [3:0] _T_585;
  wire [3:0] _T_586;
  wire  _T_588;
  wire  _T_589;
  wire  _T_591;
  wire  _T_593;
  wire [1:0] _T_594;
  wire [1:0] _T_595;
  wire  _T_596;
  wire  _T_598;
  wire  _T_600;
  wire [1:0] _T_601;
  wire [1:0] _T_602;
  wire [1:0] _T_603;
  wire [2:0] _T_604;
  wire [2:0] _T_605;
  wire [3:0] _T_606;
  wire [7:0] _T_607;
  wire [7:0] _T_608;
  wire  _T_610;
  wire [3:0] _T_611;
  wire [3:0] _T_612;
  wire  _T_614;
  wire  _T_615;
  wire  _T_617;
  wire  _T_619;
  wire [1:0] _T_620;
  wire [1:0] _T_621;
  wire  _T_622;
  wire  _T_624;
  wire  _T_626;
  wire [1:0] _T_627;
  wire [1:0] _T_628;
  wire [1:0] _T_629;
  wire [2:0] _T_630;
  wire [3:0] _T_631;
  wire [3:0] _T_632;
  wire  _T_634;
  wire  _T_635;
  wire  _T_637;
  wire  _T_639;
  wire [1:0] _T_640;
  wire [1:0] _T_641;
  wire  _T_642;
  wire  _T_644;
  wire  _T_646;
  wire [1:0] _T_647;
  wire [1:0] _T_648;
  wire [1:0] _T_649;
  wire [2:0] _T_650;
  wire [2:0] _T_651;
  wire [3:0] _T_652;
  wire [3:0] _T_653;
  wire [4:0] _T_654;
  wire [15:0] _T_655;
  wire [15:0] _T_656;
  wire  _T_658;
  wire [7:0] _T_659;
  wire [7:0] _T_660;
  wire  _T_662;
  wire [3:0] _T_663;
  wire [3:0] _T_664;
  wire  _T_666;
  wire  _T_667;
  wire  _T_669;
  wire  _T_671;
  wire [1:0] _T_672;
  wire [1:0] _T_673;
  wire  _T_674;
  wire  _T_676;
  wire  _T_678;
  wire [1:0] _T_679;
  wire [1:0] _T_680;
  wire [1:0] _T_681;
  wire [2:0] _T_682;
  wire [3:0] _T_683;
  wire [3:0] _T_684;
  wire  _T_686;
  wire  _T_687;
  wire  _T_689;
  wire  _T_691;
  wire [1:0] _T_692;
  wire [1:0] _T_693;
  wire  _T_694;
  wire  _T_696;
  wire  _T_698;
  wire [1:0] _T_699;
  wire [1:0] _T_700;
  wire [1:0] _T_701;
  wire [2:0] _T_702;
  wire [2:0] _T_703;
  wire [3:0] _T_704;
  wire [7:0] _T_705;
  wire [7:0] _T_706;
  wire  _T_708;
  wire [3:0] _T_709;
  wire [3:0] _T_710;
  wire  _T_712;
  wire  _T_713;
  wire  _T_715;
  wire  _T_717;
  wire [1:0] _T_718;
  wire [1:0] _T_719;
  wire  _T_720;
  wire  _T_722;
  wire  _T_724;
  wire [1:0] _T_725;
  wire [1:0] _T_726;
  wire [1:0] _T_727;
  wire [2:0] _T_728;
  wire [3:0] _T_729;
  wire [3:0] _T_730;
  wire  _T_732;
  wire  _T_733;
  wire  _T_735;
  wire  _T_737;
  wire [1:0] _T_738;
  wire [1:0] _T_739;
  wire  _T_740;
  wire  _T_742;
  wire  _T_744;
  wire [1:0] _T_745;
  wire [1:0] _T_746;
  wire [1:0] _T_747;
  wire [2:0] _T_748;
  wire [2:0] _T_749;
  wire [3:0] _T_750;
  wire [3:0] _T_751;
  wire [4:0] _T_752;
  wire [4:0] _T_753;
  wire [5:0] _T_754;
  wire [31:0] _T_755;
  wire [31:0] _T_756;
  wire  _T_758;
  wire [15:0] _T_759;
  wire [15:0] _T_760;
  wire  _T_762;
  wire [7:0] _T_763;
  wire [7:0] _T_764;
  wire  _T_766;
  wire [3:0] _T_767;
  wire [3:0] _T_768;
  wire  _T_770;
  wire  _T_771;
  wire  _T_773;
  wire  _T_775;
  wire [1:0] _T_776;
  wire [1:0] _T_777;
  wire  _T_778;
  wire  _T_780;
  wire  _T_782;
  wire [1:0] _T_783;
  wire [1:0] _T_784;
  wire [1:0] _T_785;
  wire [2:0] _T_786;
  wire [3:0] _T_787;
  wire [3:0] _T_788;
  wire  _T_790;
  wire  _T_791;
  wire  _T_793;
  wire  _T_795;
  wire [1:0] _T_796;
  wire [1:0] _T_797;
  wire  _T_798;
  wire  _T_800;
  wire  _T_802;
  wire [1:0] _T_803;
  wire [1:0] _T_804;
  wire [1:0] _T_805;
  wire [2:0] _T_806;
  wire [2:0] _T_807;
  wire [3:0] _T_808;
  wire [7:0] _T_809;
  wire [7:0] _T_810;
  wire  _T_812;
  wire [3:0] _T_813;
  wire [3:0] _T_814;
  wire  _T_816;
  wire  _T_817;
  wire  _T_819;
  wire  _T_821;
  wire [1:0] _T_822;
  wire [1:0] _T_823;
  wire  _T_824;
  wire  _T_826;
  wire  _T_828;
  wire [1:0] _T_829;
  wire [1:0] _T_830;
  wire [1:0] _T_831;
  wire [2:0] _T_832;
  wire [3:0] _T_833;
  wire [3:0] _T_834;
  wire  _T_836;
  wire  _T_837;
  wire  _T_839;
  wire  _T_841;
  wire [1:0] _T_842;
  wire [1:0] _T_843;
  wire  _T_844;
  wire  _T_846;
  wire  _T_848;
  wire [1:0] _T_849;
  wire [1:0] _T_850;
  wire [1:0] _T_851;
  wire [2:0] _T_852;
  wire [2:0] _T_853;
  wire [3:0] _T_854;
  wire [3:0] _T_855;
  wire [4:0] _T_856;
  wire [15:0] _T_857;
  wire [15:0] _T_858;
  wire  _T_860;
  wire [7:0] _T_861;
  wire [7:0] _T_862;
  wire  _T_864;
  wire [3:0] _T_865;
  wire [3:0] _T_866;
  wire  _T_868;
  wire  _T_869;
  wire  _T_871;
  wire  _T_873;
  wire [1:0] _T_874;
  wire [1:0] _T_875;
  wire  _T_876;
  wire  _T_878;
  wire  _T_880;
  wire [1:0] _T_881;
  wire [1:0] _T_882;
  wire [1:0] _T_883;
  wire [2:0] _T_884;
  wire [3:0] _T_885;
  wire [3:0] _T_886;
  wire  _T_888;
  wire  _T_889;
  wire  _T_891;
  wire  _T_893;
  wire [1:0] _T_894;
  wire [1:0] _T_895;
  wire  _T_896;
  wire  _T_898;
  wire  _T_900;
  wire [1:0] _T_901;
  wire [1:0] _T_902;
  wire [1:0] _T_903;
  wire [2:0] _T_904;
  wire [2:0] _T_905;
  wire [3:0] _T_906;
  wire [7:0] _T_907;
  wire [7:0] _T_908;
  wire  _T_910;
  wire [3:0] _T_911;
  wire [3:0] _T_912;
  wire  _T_914;
  wire  _T_915;
  wire  _T_917;
  wire  _T_919;
  wire [1:0] _T_920;
  wire [1:0] _T_921;
  wire  _T_922;
  wire  _T_924;
  wire  _T_926;
  wire [1:0] _T_927;
  wire [1:0] _T_928;
  wire [1:0] _T_929;
  wire [2:0] _T_930;
  wire [3:0] _T_931;
  wire [3:0] _T_932;
  wire  _T_934;
  wire  _T_935;
  wire  _T_937;
  wire  _T_939;
  wire [1:0] _T_940;
  wire [1:0] _T_941;
  wire  _T_942;
  wire  _T_944;
  wire  _T_946;
  wire [1:0] _T_947;
  wire [1:0] _T_948;
  wire [1:0] _T_949;
  wire [2:0] _T_950;
  wire [2:0] _T_951;
  wire [3:0] _T_952;
  wire [3:0] _T_953;
  wire [4:0] _T_954;
  wire [4:0] _T_955;
  wire [5:0] _T_956;
  wire [5:0] _T_957;
  wire [6:0] _T_958;
  wire [6:0] _T_959;
  wire [7:0] _T_960;
  wire [4:0] whichInterrupt;
  wire [31:0] _GEN_3;
  wire [32:0] _T_962;
  wire [31:0] interruptCause;
  wire  _T_964;
  wire  _T_965;
  wire  _T_967;
  wire  _T_968;
  wire  _T_969;
  wire [31:0] _T_971_mask;
  wire  _T_972;
  wire [30:0] _T_973;
  wire [31:0] _T_977;
  wire [30:0] _T_978;
  wire [30:0] _T_979;
  wire [30:0] _T_980;
  wire [32:0] _T_982;
  wire [31:0] _T_984_mask;
  wire  _T_985;
  wire [30:0] _T_986;
  wire [31:0] _T_990;
  wire [30:0] _T_991;
  wire [30:0] _T_992;
  wire [30:0] _T_993;
  wire [32:0] _T_995;
  wire [31:0] _T_997_mask;
  wire  _T_998;
  wire [30:0] _T_999;
  wire [31:0] _T_1003;
  wire [30:0] _T_1004;
  wire [30:0] _T_1005;
  wire [30:0] _T_1006;
  wire [32:0] _T_1008;
  wire [31:0] _T_1010_mask;
  wire  _T_1011;
  wire [30:0] _T_1012;
  wire [31:0] _T_1016;
  wire [30:0] _T_1017;
  wire [30:0] _T_1018;
  wire [30:0] _T_1019;
  wire [32:0] _T_1021;
  wire [31:0] _T_1023_mask;
  wire  _T_1024;
  wire [30:0] _T_1025;
  wire [31:0] _T_1029;
  wire [30:0] _T_1030;
  wire [30:0] _T_1031;
  wire [30:0] _T_1032;
  wire [32:0] _T_1034;
  wire [31:0] _T_1036_mask;
  wire  _T_1037;
  wire [30:0] _T_1038;
  wire [31:0] _T_1042;
  wire [30:0] _T_1043;
  wire [30:0] _T_1044;
  wire [30:0] _T_1045;
  wire [32:0] _T_1047;
  wire [31:0] _T_1049_mask;
  wire  _T_1050;
  wire [30:0] _T_1051;
  wire [31:0] _T_1055;
  wire [30:0] _T_1056;
  wire [30:0] _T_1057;
  wire [30:0] _T_1058;
  wire [32:0] _T_1060;
  wire [31:0] _T_1062_mask;
  wire  _T_1063;
  wire [30:0] _T_1064;
  wire [31:0] _T_1068;
  wire [30:0] _T_1069;
  wire [30:0] _T_1070;
  wire [30:0] _T_1071;
  wire [32:0] _T_1073;
  reg [31:0] reg_misa;
  reg [31:0] _RAND_159;
  wire [1:0] _T_1076;
  wire [2:0] _T_1077;
  wire [1:0] _T_1078;
  wire [1:0] _T_1079;
  wire [3:0] _T_1080;
  wire [6:0] _T_1081;
  wire [2:0] _T_1082;
  wire [3:0] _T_1083;
  wire [3:0] _T_1084;
  wire [2:0] _T_1085;
  wire [6:0] _T_1086;
  wire [10:0] _T_1087;
  wire [17:0] _T_1088;
  wire [1:0] _T_1089;
  wire [2:0] _T_1090;
  wire [1:0] _T_1091;
  wire [8:0] _T_1092;
  wire [10:0] _T_1093;
  wire [13:0] _T_1094;
  wire [3:0] _T_1095;
  wire [27:0] _T_1096;
  wire [31:0] _T_1097;
  wire [3:0] _T_1098;
  wire [32:0] _T_1099;
  wire [36:0] _T_1100;
  wire [68:0] _T_1101;
  wire [82:0] _T_1102;
  wire [100:0] _T_1103;
  wire [31:0] read_mstatus;
  wire [3:0] _GEN_37;
  wire  _GEN_38;
  wire [5:0] _GEN_39;
  wire [7:0] _GEN_40;
  wire  _GEN_41;
  wire  _GEN_42;
  wire [1:0] _GEN_43;
  wire [1:0] _GEN_44;
  wire  _GEN_45;
  wire  _GEN_46;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire [31:0] _GEN_52;
  wire [1:0] _T_1105;
  wire [2:0] _T_1106;
  wire [1:0] _T_1107;
  wire [1:0] _T_1108;
  wire [3:0] _T_1109;
  wire [6:0] _T_1110;
  wire [3:0] _T_1111;
  wire [1:0] _T_1112;
  wire [5:0] _T_1113;
  wire [13:0] _T_1114;
  wire [4:0] _T_1115;
  wire [18:0] _T_1116;
  wire [24:0] _T_1117;
  wire [31:0] _T_1118;
  wire [3:0] _T_1123;
  wire [5:0] _T_1124;
  wire [3:0] _T_1125;
  wire [1:0] _T_1126;
  wire [5:0] _T_1127;
  wire [11:0] _T_1128;
  wire [1:0] _T_1129;
  wire [2:0] _T_1130;
  wire [12:0] _T_1131;
  wire [3:0] _T_1132;
  wire [16:0] _T_1133;
  wire [19:0] _T_1134;
  wire [31:0] _T_1135;
  wire [31:0] _T_1139;
  wire [31:0] _T_1140;
  wire [1:0] _T_1156;
  wire [2:0] _T_1157;
  wire [2:0] _T_1158;
  wire [4:0] _T_1159;
  wire [7:0] _T_1160;
  wire [1:0] _T_1161;
  wire [2:0] _T_1162;
  wire [2:0] _T_1163;
  wire [4:0] _T_1164;
  wire [7:0] _T_1165;
  wire [1:0] _T_1166;
  wire [2:0] _T_1167;
  wire [2:0] _T_1168;
  wire [4:0] _T_1169;
  wire [7:0] _T_1170;
  wire [1:0] _T_1171;
  wire [2:0] _T_1172;
  wire [2:0] _T_1173;
  wire [4:0] _T_1174;
  wire [7:0] _T_1175;
  wire [15:0] _T_1176;
  wire [15:0] _T_1177;
  wire [31:0] _T_1178;
  wire [1:0] _T_1179;
  wire [2:0] _T_1180;
  wire [2:0] _T_1181;
  wire [4:0] _T_1182;
  wire [7:0] _T_1183;
  wire [1:0] _T_1184;
  wire [2:0] _T_1185;
  wire [2:0] _T_1186;
  wire [4:0] _T_1187;
  wire [7:0] _T_1188;
  wire [1:0] _T_1189;
  wire [2:0] _T_1190;
  wire [2:0] _T_1191;
  wire [4:0] _T_1192;
  wire [7:0] _T_1193;
  wire [1:0] _T_1194;
  wire [2:0] _T_1195;
  wire [2:0] _T_1196;
  wire [4:0] _T_1197;
  wire [7:0] _T_1198;
  wire [15:0] _T_1199;
  wire [15:0] _T_1200;
  wire [31:0] _T_1201;
  wire  _T_1249;
  wire  _T_1251;
  wire  _T_1253;
  wire  _T_1261;
  wire  _T_1263;
  wire  _T_1265;
  wire  _T_1267;
  wire  _T_1269;
  wire  _T_1271;
  wire  _T_1273;
  wire  _T_1275;
  wire  _T_1277;
  wire  _T_1279;
  wire  _T_1281;
  wire  _T_1283;
  wire  _T_1285;
  wire  _T_1287;
  wire  _T_1289;
  wire  _T_1465;
  wire  _T_1467;
  wire  _T_1469;
  wire  _T_1471;
  wire  _T_1477;
  wire  _T_1479;
  wire  _T_1481;
  wire  _T_1483;
  wire  _T_1485;
  wire  _T_1487;
  wire  _T_1489;
  wire  _T_1491;
  wire  _T_1510;
  wire  _T_1511;
  wire  _T_1512;
  wire [31:0] _T_1514;
  wire [31:0] _T_1515;
  wire [31:0] _T_1519;
  wire [31:0] _T_1520;
  wire [31:0] wdata;
  wire  system_insn;
  wire [2:0] _T_1523;
  wire [7:0] opcode;
  wire  _T_1524;
  wire  insn_call;
  wire  _T_1525;
  wire  insn_break;
  wire  _T_1526;
  wire  insn_ret;
  wire  _T_1527;
  wire  insn_wfi;
  wire [1:0] _T_1558;
  wire  _T_1559;
  wire  _T_1561;
  wire  _T_1563;
  wire  _T_1565;
  wire  _T_1567;
  wire  _T_1569;
  wire  _T_1571;
  wire  _T_1573;
  wire  _T_1575;
  wire  _T_1577;
  wire  _T_1579;
  wire  _T_1581;
  wire  _T_1583;
  wire  _T_1585;
  wire  _T_1587;
  wire  _T_1589;
  wire  _T_1591;
  wire  _T_1593;
  wire  _T_1595;
  wire  _T_1597;
  wire  _T_1599;
  wire  _T_1601;
  wire  _T_1603;
  wire  _T_1605;
  wire  _T_1607;
  wire  _T_1609;
  wire  _T_1611;
  wire  _T_1613;
  wire  _T_1615;
  wire  _T_1617;
  wire  _T_1619;
  wire  _T_1621;
  wire  _T_1623;
  wire  _T_1625;
  wire  _T_1627;
  wire  _T_1629;
  wire  _T_1631;
  wire  _T_1633;
  wire  _T_1635;
  wire  _T_1637;
  wire  _T_1639;
  wire  _T_1641;
  wire  _T_1643;
  wire  _T_1645;
  wire  _T_1647;
  wire  _T_1649;
  wire  _T_1651;
  wire  _T_1653;
  wire  _T_1655;
  wire  _T_1657;
  wire  _T_1659;
  wire  _T_1661;
  wire  _T_1663;
  wire  _T_1665;
  wire  _T_1667;
  wire  _T_1669;
  wire  _T_1671;
  wire  _T_1673;
  wire  _T_1675;
  wire  _T_1677;
  wire  _T_1679;
  wire  _T_1681;
  wire  _T_1683;
  wire  _T_1685;
  wire  _T_1687;
  wire  _T_1689;
  wire  _T_1691;
  wire  _T_1693;
  wire  _T_1695;
  wire  _T_1697;
  wire  _T_1699;
  wire  _T_1701;
  wire  _T_1703;
  wire  _T_1705;
  wire  _T_1707;
  wire  _T_1709;
  wire  _T_1711;
  wire  _T_1713;
  wire  _T_1715;
  wire  _T_1717;
  wire  _T_1719;
  wire  _T_1721;
  wire  _T_1723;
  wire  _T_1725;
  wire  _T_1727;
  wire  _T_1729;
  wire  _T_1731;
  wire  _T_1733;
  wire  _T_1735;
  wire  _T_1737;
  wire  _T_1739;
  wire  _T_1741;
  wire  _T_1743;
  wire  _T_1745;
  wire  _T_1747;
  wire  _T_1749;
  wire  _T_1751;
  wire  _T_1753;
  wire  _T_1755;
  wire  _T_1757;
  wire  _T_1759;
  wire  _T_1761;
  wire  _T_1763;
  wire  _T_1765;
  wire  _T_1767;
  wire  _T_1769;
  wire  _T_1771;
  wire  _T_1773;
  wire  _T_1775;
  wire  _T_1777;
  wire  _T_1779;
  wire  _T_1781;
  wire  _T_1783;
  wire  _T_1785;
  wire  _T_1787;
  wire  _T_1789;
  wire  _T_1791;
  wire  _T_1793;
  wire  _T_1795;
  wire  _T_1797;
  wire  _T_1799;
  wire  _T_1801;
  wire  _T_1803;
  wire  _T_1805;
  wire  _T_1807;
  wire  _T_1809;
  wire  _T_1811;
  wire  _T_1813;
  wire  _T_1815;
  wire  _T_1817;
  wire  _T_1819;
  wire  _T_1820;
  wire  _T_1821;
  wire  _T_1822;
  wire  _T_1823;
  wire  _T_1824;
  wire  _T_1825;
  wire  _T_1826;
  wire  _T_1827;
  wire  _T_1828;
  wire  _T_1829;
  wire  _T_1830;
  wire  _T_1831;
  wire  _T_1832;
  wire  _T_1833;
  wire  _T_1834;
  wire  _T_1835;
  wire  _T_1836;
  wire  _T_1837;
  wire  _T_1838;
  wire  _T_1839;
  wire  _T_1840;
  wire  _T_1841;
  wire  _T_1842;
  wire  _T_1843;
  wire  _T_1844;
  wire  _T_1845;
  wire  _T_1846;
  wire  _T_1847;
  wire  _T_1848;
  wire  _T_1849;
  wire  _T_1850;
  wire  _T_1851;
  wire  _T_1852;
  wire  _T_1853;
  wire  _T_1854;
  wire  _T_1855;
  wire  _T_1856;
  wire  _T_1857;
  wire  _T_1858;
  wire  _T_1859;
  wire  _T_1860;
  wire  _T_1861;
  wire  _T_1862;
  wire  _T_1863;
  wire  _T_1864;
  wire  _T_1865;
  wire  _T_1866;
  wire  _T_1867;
  wire  _T_1868;
  wire  _T_1869;
  wire  _T_1870;
  wire  _T_1871;
  wire  _T_1872;
  wire  _T_1873;
  wire  _T_1874;
  wire  _T_1875;
  wire  _T_1876;
  wire  _T_1877;
  wire  _T_1878;
  wire  _T_1879;
  wire  _T_1880;
  wire  _T_1881;
  wire  _T_1882;
  wire  _T_1883;
  wire  _T_1884;
  wire  _T_1885;
  wire  _T_1886;
  wire  _T_1887;
  wire  _T_1888;
  wire  _T_1889;
  wire  _T_1890;
  wire  _T_1891;
  wire  _T_1892;
  wire  _T_1893;
  wire  _T_1894;
  wire  _T_1895;
  wire  _T_1896;
  wire  _T_1897;
  wire  _T_1898;
  wire  _T_1899;
  wire  _T_1900;
  wire  _T_1901;
  wire  _T_1902;
  wire  _T_1903;
  wire  _T_1904;
  wire  _T_1905;
  wire  _T_1906;
  wire  _T_1907;
  wire  _T_1908;
  wire  _T_1909;
  wire  _T_1910;
  wire  _T_1911;
  wire  _T_1912;
  wire  _T_1913;
  wire  _T_1914;
  wire  _T_1915;
  wire  _T_1916;
  wire  _T_1917;
  wire  _T_1918;
  wire  _T_1919;
  wire  _T_1920;
  wire  _T_1921;
  wire  _T_1922;
  wire  _T_1923;
  wire  _T_1924;
  wire  _T_1925;
  wire  _T_1926;
  wire  _T_1927;
  wire  _T_1928;
  wire  _T_1929;
  wire  _T_1930;
  wire  _T_1931;
  wire  _T_1932;
  wire  _T_1933;
  wire  _T_1934;
  wire  _T_1935;
  wire  _T_1936;
  wire  _T_1937;
  wire  _T_1938;
  wire  _T_1939;
  wire  _T_1940;
  wire  _T_1941;
  wire  _T_1942;
  wire  _T_1943;
  wire  _T_1944;
  wire  _T_1945;
  wire  _T_1946;
  wire  _T_1947;
  wire  _T_1948;
  wire  _T_1950;
  wire  _T_1951;
  wire  _T_1960;
  wire  _T_1961;
  wire  _T_1962;
  wire  _T_1965;
  wire  _T_1966;
  wire  _T_1967;
  wire  _T_1968;
  wire  _T_1971;
  wire [31:0] _T_1973;
  wire  _T_1974;
  wire  _T_1975;
  wire  _T_1976;
  wire  _T_1984;
  wire  _T_1985;
  wire  _T_1989;
  wire  _T_1990;
  wire [1:0] _T_2003;
  wire [1:0] _T_2004;
  wire  _T_2006;
  wire  _T_2008;
  wire  _T_2010;
  wire  _T_2011;
  wire  _T_2013;
  wire  _T_2015;
  wire  _T_2016;
  wire  _T_2017;
  wire  _T_2019;
  wire [3:0] _GEN_4;
  wire [4:0] _T_2046;
  wire [3:0] _T_2047;
  wire [31:0] _T_2049;
  wire [31:0] cause;
  wire [4:0] cause_lsbs;
  wire  _T_2050;
  wire  _T_2052;
  wire  causeIsDebugInt;
  wire  _T_2055;
  wire  causeIsDebugTrigger;
  wire  _T_2061;
  wire [1:0] _T_2062;
  wire [1:0] _T_2063;
  wire [3:0] _T_2064;
  wire [3:0] _T_2065;
  wire  _T_2066;
  wire  causeIsDebugBreak;
  wire  _T_2068;
  wire  _T_2069;
  wire  _T_2070;
  wire  _T_2071;
  wire [11:0] _T_2074;
  wire [11:0] debugTVec;
  wire [3:0] _T_2090;
  wire [5:0] _GEN_5;
  wire [5:0] _T_2091;
  wire [25:0] _T_2092;
  wire [31:0] _T_2093;
  wire  _T_2094;
  wire  _T_2096;
  wire [31:0] notDebugTVec;
  wire [31:0] tvec;
  wire  _T_2097;
  wire  _T_2098;
  wire  _T_2101;
  wire [1:0] _T_2102;
  wire  _T_2104;
  wire [1:0] _T_2105;
  wire  _T_2107;
  wire  _T_2108;
  wire  _T_2113;
  wire [1:0] _T_2114;
  reg [1:0] _T_2116;
  reg [31:0] _RAND_160;
  wire  exception;
  wire [1:0] _T_2118;
  wire [1:0] _T_2119;
  wire [2:0] _T_2120;
  wire  _T_2122;
  wire  _T_2123;
  wire  _T_2125;
  wire  _T_2128;
  wire  _T_2131;
  wire  _GEN_53;
  wire  _T_2134;
  wire  _T_2135;
  wire  _T_2136;
  wire  _GEN_54;
  wire  _T_2139;
  wire  _T_2141;
  wire  _T_2142;
  wire  _T_2143;
  wire  _T_2145;
  wire  _T_2147;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _T_2161;
  wire  _T_2164;
  wire  _T_2165;
  wire  _T_2167;
  wire [31:0] _T_2168;
  wire [31:0] _T_2170;
  wire [31:0] _T_2171;
  wire  _T_2183;
  wire  _T_2184;
  wire  _T_2185;
  wire  _T_2186;
  wire  _T_2187;
  wire  _T_2188;
  wire  _T_2189;
  wire  _T_2190;
  wire  _T_2191;
  wire  _T_2192;
  wire  _T_2193;
  wire  _T_2194;
  wire  _T_2195;
  wire  _T_2196;
  wire  _T_2197;
  wire  _T_2198;
  wire  _T_2199;
  wire  _T_2200;
  wire  _T_2201;
  wire  _T_2202;
  wire  _T_2203;
  wire [31:0] _T_2205;
  wire [1:0] _T_2213;
  wire [1:0] _T_2214;
  wire [2:0] _T_2215;
  wire  _GEN_57;
  wire [31:0] _GEN_58;
  wire [2:0] _GEN_59;
  wire [1:0] _GEN_60;
  wire  _GEN_62;
  wire [31:0] _GEN_63;
  wire [2:0] _GEN_64;
  wire [1:0] _GEN_65;
  wire  _T_2219;
  wire [31:0] _T_2221;
  wire  _T_2222;
  wire  _T_2224;
  wire [1:0] _T_2226;
  wire [31:0] _GEN_6;
  wire [31:0] _T_2227;
  wire [31:0] _T_2228;
  wire [1:0] _GEN_71;
  wire [31:0] _GEN_74;
  wire [31:0] _GEN_75;
  wire [31:0] _GEN_76;
  wire  _GEN_77;
  wire [1:0] _GEN_78;
  wire  _GEN_79;
  wire  _GEN_81;
  wire [31:0] _GEN_82;
  wire [2:0] _GEN_83;
  wire [1:0] _GEN_84;
  wire [1:0] _GEN_90;
  wire [31:0] _GEN_92;
  wire [31:0] _GEN_93;
  wire [31:0] _GEN_94;
  wire  _GEN_95;
  wire [1:0] _GEN_96;
  wire  _GEN_97;
  wire  _T_2255;
  wire  _GEN_104;
  wire [31:0] _GEN_105;
  wire  _T_2264;
  wire  _GEN_106;
  wire  _GEN_107;
  wire [1:0] _GEN_108;
  wire [31:0] _GEN_110;
  wire [31:0] _GEN_115;
  wire  _GEN_116;
  wire  _GEN_117;
  wire  _GEN_118;
  wire [1:0] _GEN_119;
  wire  _T_2271;
  wire [31:0] _T_2273;
  wire [31:0] _T_2275;
  wire [63:0] _T_2283;
  wire [63:0] _T_2285;
  wire [31:0] _T_2287;
  wire [31:0] _T_2289;
  wire [31:0] _T_2291;
  wire [15:0] _T_2293;
  wire [31:0] _T_2295;
  wire [31:0] _T_2297;
  wire [31:0] _T_2299;
  wire [31:0] _T_2301;
  wire [31:0] _T_2303;
  wire  _T_2305;
  wire [31:0] _T_2307;
  wire [31:0] _T_2309;
  wire [31:0] _T_2311;
  wire [31:0] _T_2487;
  wire [31:0] _T_2489;
  wire [31:0] _T_2491;
  wire [31:0] _T_2493;
  wire [29:0] _T_2499;
  wire [29:0] _T_2501;
  wire [29:0] _T_2503;
  wire [29:0] _T_2505;
  wire [29:0] _T_2507;
  wire [29:0] _T_2509;
  wire [29:0] _T_2511;
  wire [29:0] _T_2513;
  wire [31:0] _GEN_8;
  wire [31:0] _T_2530;
  wire [31:0] _T_2531;
  wire [63:0] _GEN_9;
  wire [63:0] _T_2535;
  wire [63:0] _T_2536;
  wire [63:0] _GEN_10;
  wire [63:0] _T_2537;
  wire [63:0] _GEN_11;
  wire [63:0] _T_2538;
  wire [63:0] _GEN_12;
  wire [63:0] _T_2539;
  wire [63:0] _GEN_13;
  wire [63:0] _T_2540;
  wire [63:0] _GEN_14;
  wire [63:0] _T_2541;
  wire [63:0] _GEN_15;
  wire [63:0] _T_2542;
  wire [63:0] _GEN_16;
  wire [63:0] _T_2543;
  wire [63:0] _GEN_431;
  wire [63:0] _T_2544;
  wire [63:0] _GEN_432;
  wire [63:0] _T_2545;
  wire [63:0] _GEN_433;
  wire [63:0] _T_2546;
  wire [63:0] _GEN_434;
  wire [63:0] _T_2547;
  wire [63:0] _GEN_435;
  wire [63:0] _T_2548;
  wire [63:0] _GEN_436;
  wire [63:0] _T_2549;
  wire [63:0] _GEN_437;
  wire [63:0] _T_2637;
  wire [63:0] _GEN_438;
  wire [63:0] _T_2638;
  wire [63:0] _GEN_439;
  wire [63:0] _T_2639;
  wire [63:0] _GEN_440;
  wire [63:0] _T_2640;
  wire [63:0] _GEN_441;
  wire [63:0] _T_2643;
  wire [63:0] _GEN_442;
  wire [63:0] _T_2644;
  wire [63:0] _GEN_443;
  wire [63:0] _T_2645;
  wire [63:0] _GEN_444;
  wire [63:0] _T_2646;
  wire [63:0] _GEN_445;
  wire [63:0] _T_2647;
  wire [63:0] _GEN_446;
  wire [63:0] _T_2648;
  wire [63:0] _GEN_447;
  wire [63:0] _T_2649;
  wire [63:0] _GEN_448;
  wire [63:0] _T_2650;
  wire  _T_2667;
  wire  _T_2669;
  wire [100:0] _T_2674;
  wire  _T_2678;
  wire  _T_2682;
  wire  _GEN_121;
  wire  _GEN_122;
  wire  _T_2705;
  wire [31:0] _T_2706;
  wire  _T_2708;
  wire [3:0] _GEN_449;
  wire [3:0] _T_2709;
  wire [31:0] _GEN_450;
  wire [31:0] _T_2710;
  wire [31:0] _T_2711;
  wire [31:0] _T_2712;
  wire [31:0] _T_2714;
  wire [31:0] _T_2715;
  wire [31:0] _GEN_123;
  wire [31:0] _T_2772;
  wire [31:0] _GEN_124;
  wire [31:0] _T_2779;
  wire [31:0] _T_2780;
  wire [31:0] _GEN_125;
  wire [31:0] _GEN_126;
  wire [31:0] _T_2783;
  wire  _T_2784;
  wire [5:0] _T_2787;
  wire [31:0] _GEN_453;
  wire [31:0] _T_2788;
  wire [31:0] _T_2789;
  wire [31:0] _GEN_127;
  wire [31:0] _T_2791;
  wire [31:0] _GEN_128;
  wire [31:0] _GEN_129;
  wire [31:0] _T_2793;
  wire [63:0] _T_2794;
  wire [57:0] _T_2795;
  wire [63:0] _GEN_130;
  wire [57:0] _GEN_131;
  wire [31:0] _T_2797;
  wire [63:0] _T_2798;
  wire [57:0] _T_2799;
  wire [63:0] _GEN_132;
  wire [57:0] _GEN_133;
  wire [31:0] _T_2800;
  wire [63:0] _T_2801;
  wire [57:0] _T_2802;
  wire [63:0] _GEN_134;
  wire [57:0] _GEN_135;
  wire [31:0] _T_2804;
  wire [63:0] _T_2805;
  wire [57:0] _T_2806;
  wire [63:0] _GEN_136;
  wire [57:0] _GEN_137;
  wire  _T_2813;
  wire  _T_2819;
  wire  _T_2822;
  wire  _GEN_138;
  wire  _GEN_139;
  wire [31:0] _T_2828;
  wire [31:0] _T_2829;
  wire [31:0] _GEN_140;
  wire [31:0] _GEN_141;
  wire  _T_2832;
  wire  _T_2833;
  wire  _T_2840;
  wire [1:0] _T_2846;
  wire  _T_2852;
  wire  _T_2854;
  wire  _GEN_145;
  wire  _GEN_151;
  wire [1:0] _GEN_157;
  wire  _GEN_167;
  wire  _GEN_169;
  wire  _GEN_171;
  wire  _GEN_173;
  wire  _T_2855;
  wire  _GEN_175;
  wire  _GEN_179;
  wire  _GEN_185;
  wire [1:0] _GEN_191;
  wire  _GEN_201;
  wire  _GEN_203;
  wire  _GEN_205;
  wire [31:0] _GEN_207;
  wire [31:0] _GEN_209;
  wire  _GEN_213;
  wire  _GEN_219;
  wire [1:0] _GEN_225;
  wire  _GEN_235;
  wire  _GEN_237;
  wire  _GEN_239;
  wire [31:0] _GEN_241;
  wire  _T_2857;
  wire  _T_2858;
  wire [7:0] _T_2864;
  wire  _T_2865;
  wire  _T_2866;
  wire  _T_2867;
  wire [1:0] _T_2868;
  wire  _T_2870;
  wire  _GEN_243;
  wire [1:0] _GEN_245;
  wire  _GEN_246;
  wire  _GEN_247;
  wire  _GEN_248;
  wire  _T_2871;
  wire  _T_2872;
  wire  _T_2873;
  wire  _T_2875;
  wire  _T_2876;
  wire [31:0] _GEN_249;
  wire  _T_2878;
  wire  _T_2879;
  wire [23:0] _T_2881;
  wire [7:0] _T_2885;
  wire  _T_2886;
  wire  _T_2887;
  wire  _T_2888;
  wire [1:0] _T_2889;
  wire  _T_2891;
  wire  _GEN_250;
  wire [1:0] _GEN_252;
  wire  _GEN_253;
  wire  _GEN_254;
  wire  _GEN_255;
  wire  _T_2892;
  wire  _T_2893;
  wire  _T_2894;
  wire  _T_2896;
  wire  _T_2897;
  wire [31:0] _GEN_256;
  wire  _T_2899;
  wire  _T_2900;
  wire [15:0] _T_2902;
  wire [7:0] _T_2906;
  wire  _T_2907;
  wire  _T_2908;
  wire  _T_2909;
  wire [1:0] _T_2910;
  wire  _T_2912;
  wire  _GEN_257;
  wire [1:0] _GEN_259;
  wire  _GEN_260;
  wire  _GEN_261;
  wire  _GEN_262;
  wire  _T_2913;
  wire  _T_2914;
  wire  _T_2915;
  wire  _T_2917;
  wire  _T_2918;
  wire [31:0] _GEN_263;
  wire  _T_2920;
  wire  _T_2921;
  wire [7:0] _T_2923;
  wire  _T_2928;
  wire  _T_2929;
  wire  _T_2930;
  wire [1:0] _T_2931;
  wire  _T_2933;
  wire  _GEN_264;
  wire [1:0] _GEN_266;
  wire  _GEN_267;
  wire  _GEN_268;
  wire  _GEN_269;
  wire  _T_2934;
  wire  _T_2935;
  wire  _T_2936;
  wire  _T_2938;
  wire  _T_2939;
  wire [31:0] _GEN_270;
  wire  _T_2941;
  wire  _T_2942;
  wire [7:0] _T_2948;
  wire  _T_2949;
  wire  _T_2950;
  wire  _T_2951;
  wire [1:0] _T_2952;
  wire  _T_2954;
  wire  _GEN_271;
  wire [1:0] _GEN_273;
  wire  _GEN_274;
  wire  _GEN_275;
  wire  _GEN_276;
  wire  _T_2955;
  wire  _T_2956;
  wire  _T_2957;
  wire  _T_2959;
  wire  _T_2960;
  wire [31:0] _GEN_277;
  wire  _T_2962;
  wire  _T_2963;
  wire [7:0] _T_2969;
  wire  _T_2970;
  wire  _T_2971;
  wire  _T_2972;
  wire [1:0] _T_2973;
  wire  _T_2975;
  wire  _GEN_278;
  wire [1:0] _GEN_280;
  wire  _GEN_281;
  wire  _GEN_282;
  wire  _GEN_283;
  wire  _T_2976;
  wire  _T_2977;
  wire  _T_2978;
  wire  _T_2980;
  wire  _T_2981;
  wire [31:0] _GEN_284;
  wire  _T_2983;
  wire  _T_2984;
  wire [7:0] _T_2990;
  wire  _T_2991;
  wire  _T_2992;
  wire  _T_2993;
  wire [1:0] _T_2994;
  wire  _T_2996;
  wire  _GEN_285;
  wire [1:0] _GEN_287;
  wire  _GEN_288;
  wire  _GEN_289;
  wire  _GEN_290;
  wire  _T_2997;
  wire  _T_2998;
  wire  _T_2999;
  wire  _T_3001;
  wire  _T_3002;
  wire [31:0] _GEN_291;
  wire  _T_3004;
  wire  _T_3005;
  wire  _GEN_292;
  wire [1:0] _GEN_294;
  wire  _GEN_295;
  wire  _GEN_296;
  wire  _GEN_297;
  wire  _T_3020;
  wire  _T_3022;
  wire  _T_3023;
  wire [31:0] _GEN_298;
  wire  _GEN_299;
  wire  _GEN_300;
  wire [31:0] _GEN_301;
  wire [31:0] _GEN_302;
  wire [31:0] _GEN_303;
  wire [31:0] _GEN_304;
  wire [31:0] _GEN_305;
  wire [31:0] _GEN_306;
  wire [31:0] _GEN_307;
  wire [63:0] _GEN_308;
  wire [57:0] _GEN_309;
  wire [63:0] _GEN_310;
  wire [57:0] _GEN_311;
  wire  _GEN_312;
  wire  _GEN_313;
  wire [31:0] _GEN_314;
  wire [31:0] _GEN_315;
  wire  _GEN_319;
  wire  _GEN_325;
  wire [1:0] _GEN_331;
  wire  _GEN_341;
  wire  _GEN_343;
  wire  _GEN_345;
  wire [31:0] _GEN_347;
  wire  _GEN_349;
  wire [1:0] _GEN_351;
  wire  _GEN_352;
  wire  _GEN_353;
  wire  _GEN_354;
  wire [31:0] _GEN_355;
  wire  _GEN_356;
  wire [1:0] _GEN_358;
  wire  _GEN_359;
  wire  _GEN_360;
  wire  _GEN_361;
  wire [31:0] _GEN_362;
  wire  _GEN_363;
  wire [1:0] _GEN_365;
  wire  _GEN_366;
  wire  _GEN_367;
  wire  _GEN_368;
  wire [31:0] _GEN_369;
  wire  _GEN_370;
  wire [1:0] _GEN_372;
  wire  _GEN_373;
  wire  _GEN_374;
  wire  _GEN_375;
  wire [31:0] _GEN_376;
  wire  _GEN_377;
  wire [1:0] _GEN_379;
  wire  _GEN_380;
  wire  _GEN_381;
  wire  _GEN_382;
  wire [31:0] _GEN_383;
  wire  _GEN_384;
  wire [1:0] _GEN_386;
  wire  _GEN_387;
  wire  _GEN_388;
  wire  _GEN_389;
  wire [31:0] _GEN_390;
  wire  _GEN_391;
  wire [1:0] _GEN_393;
  wire  _GEN_394;
  wire  _GEN_395;
  wire  _GEN_396;
  wire [31:0] _GEN_397;
  wire  _GEN_398;
  wire [1:0] _GEN_400;
  wire  _GEN_401;
  wire  _GEN_402;
  wire  _GEN_403;
  wire [31:0] _GEN_404;
  wire  _GEN_405;
  wire  _GEN_406;
  wire  _GEN_407;
  wire  _GEN_408;
  wire  _GEN_409;
  wire [1:0] _GEN_415;
  wire  _GEN_416;
  wire [1:0] _GEN_417;
  wire  _GEN_418;
  wire [1:0] _GEN_419;
  wire  _GEN_420;
  wire [1:0] _GEN_421;
  wire  _GEN_422;
  wire [1:0] _GEN_423;
  wire  _GEN_424;
  wire [1:0] _GEN_425;
  wire  _GEN_426;
  wire [1:0] _GEN_427;
  wire  _GEN_428;
  wire [1:0] _GEN_429;
  wire  _GEN_430;
  assign io_rw_rdata = _T_2650[31:0];
  assign io_decode_read_illegal = _T_1990;
  assign io_decode_write_illegal = _T_2006;
  assign io_decode_write_flush = _T_2019;
  assign io_decode_system_illegal = _T_1559;
  assign io_csr_stall = reg_wfi;
  assign io_eret = _T_2098;
  assign io_singleStep = _T_2101;
  assign io_status_debug = reg_debug;
  assign io_status_isa = reg_misa;
  assign io_status_dprv = _T_2116;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = _T_2108;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign io_status_sxl = 2'h0;
  assign io_status_uxl = 2'h0;
  assign io_status_sd_rv32 = io_status_sd;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign io_status_tsr = reg_mstatus_tsr;
  assign io_status_tw = reg_mstatus_tw;
  assign io_status_tvm = reg_mstatus_tvm;
  assign io_status_mxr = reg_mstatus_mxr;
  assign io_status_sum = reg_mstatus_sum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = reg_mstatus_xs;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = reg_mstatus_hpp;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = reg_mstatus_hpie;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = reg_mstatus_upie;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = reg_mstatus_hie;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = reg_mstatus_uie;
  assign io_ptbr_ppn = reg_sptbr_ppn;
  assign io_evec = _GEN_115;
  assign io_time = _T_270[31:0];
  assign io_interrupt = _T_969;
  assign io_interrupt_cause = interruptCause;
  assign io_bp_0_control_action = reg_bp_0_control_action;
  assign io_bp_0_control_chain = reg_bp_0_control_chain;
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_h = reg_bp_0_control_h;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_address = reg_bp_0_address;
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l;
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a;
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x;
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w;
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r;
  assign io_pmp_0_addr = reg_pmp_0_addr;
  assign io_pmp_0_mask = _T_971_mask;
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l;
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a;
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x;
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w;
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r;
  assign io_pmp_1_addr = reg_pmp_1_addr;
  assign io_pmp_1_mask = _T_984_mask;
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l;
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a;
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x;
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w;
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r;
  assign io_pmp_2_addr = reg_pmp_2_addr;
  assign io_pmp_2_mask = _T_997_mask;
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l;
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a;
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x;
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w;
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r;
  assign io_pmp_3_addr = reg_pmp_3_addr;
  assign io_pmp_3_mask = _T_1010_mask;
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l;
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a;
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x;
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w;
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r;
  assign io_pmp_4_addr = reg_pmp_4_addr;
  assign io_pmp_4_mask = _T_1023_mask;
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l;
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a;
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x;
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w;
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r;
  assign io_pmp_5_addr = reg_pmp_5_addr;
  assign io_pmp_5_mask = _T_1036_mask;
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l;
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a;
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x;
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w;
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r;
  assign io_pmp_6_addr = reg_pmp_6_addr;
  assign io_pmp_6_mask = _T_1049_mask;
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l;
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a;
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x;
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w;
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r;
  assign io_pmp_7_addr = reg_pmp_7_addr;
  assign io_pmp_7_mask = _T_1062_mask;
  assign _GEN_0 = {{5'd0}, io_retire};
  assign _T_249 = _T_248 + _GEN_0;
  assign _T_253 = _T_249[6];
  assign _T_255 = _T_252 + 58'h1;
  assign _T_256 = _T_255[57:0];
  assign _GEN_35 = _T_253 ? _T_256 : _T_252;
  assign _T_257 = {_T_252,_T_248};
  assign _T_262 = _T_261 + 6'h1;
  assign _T_266 = _T_262[6];
  assign _T_268 = _T_265 + 58'h1;
  assign _T_269 = _T_268[57:0];
  assign _GEN_36 = _T_266 ? _T_269 : _T_265;
  assign _T_270 = {_T_265,_T_261};
  assign _T_273 = reg_mstatus_prv == 2'h1;
  assign hpm_mask = reg_mcounteren & 32'h7;
  assign _T_282 = {reg_mip_ssip,reg_mip_usip};
  assign _T_283 = {reg_mip_msip,reg_mip_hsip};
  assign _T_284 = {_T_283,_T_282};
  assign _T_285 = {reg_mip_stip,reg_mip_utip};
  assign _T_286 = {reg_mip_mtip,reg_mip_htip};
  assign _T_287 = {_T_286,_T_285};
  assign _T_288 = {_T_287,_T_284};
  assign _T_289 = {reg_mip_seip,reg_mip_ueip};
  assign _T_290 = {reg_mip_meip,reg_mip_heip};
  assign _T_291 = {_T_290,_T_289};
  assign _T_292 = {reg_mip_zero1,io_rocc_interrupt};
  assign _T_293 = {reg_mip_zero2,reg_mip_debug};
  assign _T_294 = {_T_293,_T_292};
  assign _T_295 = {_T_294,_T_291};
  assign _T_296 = {_T_295,_T_288};
  assign read_mip = _T_296 & 16'h888;
  assign _GEN_1 = {{16'd0}, read_mip};
  assign pending_interrupts = _GEN_1 & reg_mie;
  assign _GEN_2 = {{14'd0}, reg_debugint};
  assign d_interrupts = _GEN_2 << 14;
  assign _T_298 = reg_mstatus_prv <= 2'h1;
  assign _T_300 = reg_mstatus_prv == 2'h3;
  assign _T_301 = _T_300 & reg_mstatus_mie;
  assign _T_302 = _T_298 | _T_301;
  assign _T_303 = ~ reg_mideleg;
  assign _T_304 = pending_interrupts & _T_303;
  assign m_interrupts = _T_302 ? _T_304 : 32'h0;
  assign _T_307 = m_interrupts == 32'h0;
  assign _T_309 = reg_mstatus_prv < 2'h1;
  assign _T_312 = _T_273 & reg_mstatus_sie;
  assign _T_313 = _T_309 | _T_312;
  assign _T_314 = _T_307 & _T_313;
  assign _T_315 = pending_interrupts & reg_mideleg;
  assign s_interrupts = _T_314 ? _T_315 : 32'h0;
  assign _T_319 = s_interrupts & 32'hffffff0f;
  assign _T_320 = s_interrupts & 32'hf0;
  assign _T_321 = {_T_319,_T_320};
  assign _T_323 = m_interrupts & 32'hffffff0f;
  assign _T_324 = m_interrupts & 32'hf0;
  assign _T_325 = {_T_323,_T_324};
  assign _T_327 = {17'h0,d_interrupts};
  assign _T_329 = _T_327 & 32'hffffff0f;
  assign _T_332 = _T_327 & 32'hf0;
  assign _T_333 = {_T_329,_T_332};
  assign _T_335 = s_interrupts != 32'h0;
  assign _T_337 = m_interrupts != 32'h0;
  assign _T_339 = d_interrupts != 15'h0;
  assign _T_340 = _T_335 | _T_337;
  assign anyInterrupt = _T_340 | _T_339;
  assign _T_341 = {_T_333,_T_325};
  assign _T_342 = {_T_341,_T_321};
  assign _T_343 = _T_342[191:128];
  assign _T_344 = _T_342[127:0];
  assign _T_346 = _T_343 != 64'h0;
  assign _T_347 = _T_343[63:32];
  assign _T_348 = _T_343[31:0];
  assign _T_350 = _T_347 != 32'h0;
  assign _T_351 = _T_347[31:16];
  assign _T_352 = _T_347[15:0];
  assign _T_354 = _T_351 != 16'h0;
  assign _T_355 = _T_351[15:8];
  assign _T_356 = _T_351[7:0];
  assign _T_358 = _T_355 != 8'h0;
  assign _T_359 = _T_355[7:4];
  assign _T_360 = _T_355[3:0];
  assign _T_362 = _T_359 != 4'h0;
  assign _T_363 = _T_359[3];
  assign _T_365 = _T_359[2];
  assign _T_367 = _T_359[1];
  assign _T_368 = _T_365 ? 2'h2 : {{1'd0}, _T_367};
  assign _T_369 = _T_363 ? 2'h3 : _T_368;
  assign _T_370 = _T_360[3];
  assign _T_372 = _T_360[2];
  assign _T_374 = _T_360[1];
  assign _T_375 = _T_372 ? 2'h2 : {{1'd0}, _T_374};
  assign _T_376 = _T_370 ? 2'h3 : _T_375;
  assign _T_377 = _T_362 ? _T_369 : _T_376;
  assign _T_378 = {_T_362,_T_377};
  assign _T_379 = _T_356[7:4];
  assign _T_380 = _T_356[3:0];
  assign _T_382 = _T_379 != 4'h0;
  assign _T_383 = _T_379[3];
  assign _T_385 = _T_379[2];
  assign _T_387 = _T_379[1];
  assign _T_388 = _T_385 ? 2'h2 : {{1'd0}, _T_387};
  assign _T_389 = _T_383 ? 2'h3 : _T_388;
  assign _T_390 = _T_380[3];
  assign _T_392 = _T_380[2];
  assign _T_394 = _T_380[1];
  assign _T_395 = _T_392 ? 2'h2 : {{1'd0}, _T_394};
  assign _T_396 = _T_390 ? 2'h3 : _T_395;
  assign _T_397 = _T_382 ? _T_389 : _T_396;
  assign _T_398 = {_T_382,_T_397};
  assign _T_399 = _T_358 ? _T_378 : _T_398;
  assign _T_400 = {_T_358,_T_399};
  assign _T_401 = _T_352[15:8];
  assign _T_402 = _T_352[7:0];
  assign _T_404 = _T_401 != 8'h0;
  assign _T_405 = _T_401[7:4];
  assign _T_406 = _T_401[3:0];
  assign _T_408 = _T_405 != 4'h0;
  assign _T_409 = _T_405[3];
  assign _T_411 = _T_405[2];
  assign _T_413 = _T_405[1];
  assign _T_414 = _T_411 ? 2'h2 : {{1'd0}, _T_413};
  assign _T_415 = _T_409 ? 2'h3 : _T_414;
  assign _T_416 = _T_406[3];
  assign _T_418 = _T_406[2];
  assign _T_420 = _T_406[1];
  assign _T_421 = _T_418 ? 2'h2 : {{1'd0}, _T_420};
  assign _T_422 = _T_416 ? 2'h3 : _T_421;
  assign _T_423 = _T_408 ? _T_415 : _T_422;
  assign _T_424 = {_T_408,_T_423};
  assign _T_425 = _T_402[7:4];
  assign _T_426 = _T_402[3:0];
  assign _T_428 = _T_425 != 4'h0;
  assign _T_429 = _T_425[3];
  assign _T_431 = _T_425[2];
  assign _T_433 = _T_425[1];
  assign _T_434 = _T_431 ? 2'h2 : {{1'd0}, _T_433};
  assign _T_435 = _T_429 ? 2'h3 : _T_434;
  assign _T_436 = _T_426[3];
  assign _T_438 = _T_426[2];
  assign _T_440 = _T_426[1];
  assign _T_441 = _T_438 ? 2'h2 : {{1'd0}, _T_440};
  assign _T_442 = _T_436 ? 2'h3 : _T_441;
  assign _T_443 = _T_428 ? _T_435 : _T_442;
  assign _T_444 = {_T_428,_T_443};
  assign _T_445 = _T_404 ? _T_424 : _T_444;
  assign _T_446 = {_T_404,_T_445};
  assign _T_447 = _T_354 ? _T_400 : _T_446;
  assign _T_448 = {_T_354,_T_447};
  assign _T_449 = _T_348[31:16];
  assign _T_450 = _T_348[15:0];
  assign _T_452 = _T_449 != 16'h0;
  assign _T_453 = _T_449[15:8];
  assign _T_454 = _T_449[7:0];
  assign _T_456 = _T_453 != 8'h0;
  assign _T_457 = _T_453[7:4];
  assign _T_458 = _T_453[3:0];
  assign _T_460 = _T_457 != 4'h0;
  assign _T_461 = _T_457[3];
  assign _T_463 = _T_457[2];
  assign _T_465 = _T_457[1];
  assign _T_466 = _T_463 ? 2'h2 : {{1'd0}, _T_465};
  assign _T_467 = _T_461 ? 2'h3 : _T_466;
  assign _T_468 = _T_458[3];
  assign _T_470 = _T_458[2];
  assign _T_472 = _T_458[1];
  assign _T_473 = _T_470 ? 2'h2 : {{1'd0}, _T_472};
  assign _T_474 = _T_468 ? 2'h3 : _T_473;
  assign _T_475 = _T_460 ? _T_467 : _T_474;
  assign _T_476 = {_T_460,_T_475};
  assign _T_477 = _T_454[7:4];
  assign _T_478 = _T_454[3:0];
  assign _T_480 = _T_477 != 4'h0;
  assign _T_481 = _T_477[3];
  assign _T_483 = _T_477[2];
  assign _T_485 = _T_477[1];
  assign _T_486 = _T_483 ? 2'h2 : {{1'd0}, _T_485};
  assign _T_487 = _T_481 ? 2'h3 : _T_486;
  assign _T_488 = _T_478[3];
  assign _T_490 = _T_478[2];
  assign _T_492 = _T_478[1];
  assign _T_493 = _T_490 ? 2'h2 : {{1'd0}, _T_492};
  assign _T_494 = _T_488 ? 2'h3 : _T_493;
  assign _T_495 = _T_480 ? _T_487 : _T_494;
  assign _T_496 = {_T_480,_T_495};
  assign _T_497 = _T_456 ? _T_476 : _T_496;
  assign _T_498 = {_T_456,_T_497};
  assign _T_499 = _T_450[15:8];
  assign _T_500 = _T_450[7:0];
  assign _T_502 = _T_499 != 8'h0;
  assign _T_503 = _T_499[7:4];
  assign _T_504 = _T_499[3:0];
  assign _T_506 = _T_503 != 4'h0;
  assign _T_507 = _T_503[3];
  assign _T_509 = _T_503[2];
  assign _T_511 = _T_503[1];
  assign _T_512 = _T_509 ? 2'h2 : {{1'd0}, _T_511};
  assign _T_513 = _T_507 ? 2'h3 : _T_512;
  assign _T_514 = _T_504[3];
  assign _T_516 = _T_504[2];
  assign _T_518 = _T_504[1];
  assign _T_519 = _T_516 ? 2'h2 : {{1'd0}, _T_518};
  assign _T_520 = _T_514 ? 2'h3 : _T_519;
  assign _T_521 = _T_506 ? _T_513 : _T_520;
  assign _T_522 = {_T_506,_T_521};
  assign _T_523 = _T_500[7:4];
  assign _T_524 = _T_500[3:0];
  assign _T_526 = _T_523 != 4'h0;
  assign _T_527 = _T_523[3];
  assign _T_529 = _T_523[2];
  assign _T_531 = _T_523[1];
  assign _T_532 = _T_529 ? 2'h2 : {{1'd0}, _T_531};
  assign _T_533 = _T_527 ? 2'h3 : _T_532;
  assign _T_534 = _T_524[3];
  assign _T_536 = _T_524[2];
  assign _T_538 = _T_524[1];
  assign _T_539 = _T_536 ? 2'h2 : {{1'd0}, _T_538};
  assign _T_540 = _T_534 ? 2'h3 : _T_539;
  assign _T_541 = _T_526 ? _T_533 : _T_540;
  assign _T_542 = {_T_526,_T_541};
  assign _T_543 = _T_502 ? _T_522 : _T_542;
  assign _T_544 = {_T_502,_T_543};
  assign _T_545 = _T_452 ? _T_498 : _T_544;
  assign _T_546 = {_T_452,_T_545};
  assign _T_547 = _T_350 ? _T_448 : _T_546;
  assign _T_548 = {_T_350,_T_547};
  assign _T_549 = _T_344[127:64];
  assign _T_550 = _T_344[63:0];
  assign _T_552 = _T_549 != 64'h0;
  assign _T_553 = _T_549[63:32];
  assign _T_554 = _T_549[31:0];
  assign _T_556 = _T_553 != 32'h0;
  assign _T_557 = _T_553[31:16];
  assign _T_558 = _T_553[15:0];
  assign _T_560 = _T_557 != 16'h0;
  assign _T_561 = _T_557[15:8];
  assign _T_562 = _T_557[7:0];
  assign _T_564 = _T_561 != 8'h0;
  assign _T_565 = _T_561[7:4];
  assign _T_566 = _T_561[3:0];
  assign _T_568 = _T_565 != 4'h0;
  assign _T_569 = _T_565[3];
  assign _T_571 = _T_565[2];
  assign _T_573 = _T_565[1];
  assign _T_574 = _T_571 ? 2'h2 : {{1'd0}, _T_573};
  assign _T_575 = _T_569 ? 2'h3 : _T_574;
  assign _T_576 = _T_566[3];
  assign _T_578 = _T_566[2];
  assign _T_580 = _T_566[1];
  assign _T_581 = _T_578 ? 2'h2 : {{1'd0}, _T_580};
  assign _T_582 = _T_576 ? 2'h3 : _T_581;
  assign _T_583 = _T_568 ? _T_575 : _T_582;
  assign _T_584 = {_T_568,_T_583};
  assign _T_585 = _T_562[7:4];
  assign _T_586 = _T_562[3:0];
  assign _T_588 = _T_585 != 4'h0;
  assign _T_589 = _T_585[3];
  assign _T_591 = _T_585[2];
  assign _T_593 = _T_585[1];
  assign _T_594 = _T_591 ? 2'h2 : {{1'd0}, _T_593};
  assign _T_595 = _T_589 ? 2'h3 : _T_594;
  assign _T_596 = _T_586[3];
  assign _T_598 = _T_586[2];
  assign _T_600 = _T_586[1];
  assign _T_601 = _T_598 ? 2'h2 : {{1'd0}, _T_600};
  assign _T_602 = _T_596 ? 2'h3 : _T_601;
  assign _T_603 = _T_588 ? _T_595 : _T_602;
  assign _T_604 = {_T_588,_T_603};
  assign _T_605 = _T_564 ? _T_584 : _T_604;
  assign _T_606 = {_T_564,_T_605};
  assign _T_607 = _T_558[15:8];
  assign _T_608 = _T_558[7:0];
  assign _T_610 = _T_607 != 8'h0;
  assign _T_611 = _T_607[7:4];
  assign _T_612 = _T_607[3:0];
  assign _T_614 = _T_611 != 4'h0;
  assign _T_615 = _T_611[3];
  assign _T_617 = _T_611[2];
  assign _T_619 = _T_611[1];
  assign _T_620 = _T_617 ? 2'h2 : {{1'd0}, _T_619};
  assign _T_621 = _T_615 ? 2'h3 : _T_620;
  assign _T_622 = _T_612[3];
  assign _T_624 = _T_612[2];
  assign _T_626 = _T_612[1];
  assign _T_627 = _T_624 ? 2'h2 : {{1'd0}, _T_626};
  assign _T_628 = _T_622 ? 2'h3 : _T_627;
  assign _T_629 = _T_614 ? _T_621 : _T_628;
  assign _T_630 = {_T_614,_T_629};
  assign _T_631 = _T_608[7:4];
  assign _T_632 = _T_608[3:0];
  assign _T_634 = _T_631 != 4'h0;
  assign _T_635 = _T_631[3];
  assign _T_637 = _T_631[2];
  assign _T_639 = _T_631[1];
  assign _T_640 = _T_637 ? 2'h2 : {{1'd0}, _T_639};
  assign _T_641 = _T_635 ? 2'h3 : _T_640;
  assign _T_642 = _T_632[3];
  assign _T_644 = _T_632[2];
  assign _T_646 = _T_632[1];
  assign _T_647 = _T_644 ? 2'h2 : {{1'd0}, _T_646};
  assign _T_648 = _T_642 ? 2'h3 : _T_647;
  assign _T_649 = _T_634 ? _T_641 : _T_648;
  assign _T_650 = {_T_634,_T_649};
  assign _T_651 = _T_610 ? _T_630 : _T_650;
  assign _T_652 = {_T_610,_T_651};
  assign _T_653 = _T_560 ? _T_606 : _T_652;
  assign _T_654 = {_T_560,_T_653};
  assign _T_655 = _T_554[31:16];
  assign _T_656 = _T_554[15:0];
  assign _T_658 = _T_655 != 16'h0;
  assign _T_659 = _T_655[15:8];
  assign _T_660 = _T_655[7:0];
  assign _T_662 = _T_659 != 8'h0;
  assign _T_663 = _T_659[7:4];
  assign _T_664 = _T_659[3:0];
  assign _T_666 = _T_663 != 4'h0;
  assign _T_667 = _T_663[3];
  assign _T_669 = _T_663[2];
  assign _T_671 = _T_663[1];
  assign _T_672 = _T_669 ? 2'h2 : {{1'd0}, _T_671};
  assign _T_673 = _T_667 ? 2'h3 : _T_672;
  assign _T_674 = _T_664[3];
  assign _T_676 = _T_664[2];
  assign _T_678 = _T_664[1];
  assign _T_679 = _T_676 ? 2'h2 : {{1'd0}, _T_678};
  assign _T_680 = _T_674 ? 2'h3 : _T_679;
  assign _T_681 = _T_666 ? _T_673 : _T_680;
  assign _T_682 = {_T_666,_T_681};
  assign _T_683 = _T_660[7:4];
  assign _T_684 = _T_660[3:0];
  assign _T_686 = _T_683 != 4'h0;
  assign _T_687 = _T_683[3];
  assign _T_689 = _T_683[2];
  assign _T_691 = _T_683[1];
  assign _T_692 = _T_689 ? 2'h2 : {{1'd0}, _T_691};
  assign _T_693 = _T_687 ? 2'h3 : _T_692;
  assign _T_694 = _T_684[3];
  assign _T_696 = _T_684[2];
  assign _T_698 = _T_684[1];
  assign _T_699 = _T_696 ? 2'h2 : {{1'd0}, _T_698};
  assign _T_700 = _T_694 ? 2'h3 : _T_699;
  assign _T_701 = _T_686 ? _T_693 : _T_700;
  assign _T_702 = {_T_686,_T_701};
  assign _T_703 = _T_662 ? _T_682 : _T_702;
  assign _T_704 = {_T_662,_T_703};
  assign _T_705 = _T_656[15:8];
  assign _T_706 = _T_656[7:0];
  assign _T_708 = _T_705 != 8'h0;
  assign _T_709 = _T_705[7:4];
  assign _T_710 = _T_705[3:0];
  assign _T_712 = _T_709 != 4'h0;
  assign _T_713 = _T_709[3];
  assign _T_715 = _T_709[2];
  assign _T_717 = _T_709[1];
  assign _T_718 = _T_715 ? 2'h2 : {{1'd0}, _T_717};
  assign _T_719 = _T_713 ? 2'h3 : _T_718;
  assign _T_720 = _T_710[3];
  assign _T_722 = _T_710[2];
  assign _T_724 = _T_710[1];
  assign _T_725 = _T_722 ? 2'h2 : {{1'd0}, _T_724};
  assign _T_726 = _T_720 ? 2'h3 : _T_725;
  assign _T_727 = _T_712 ? _T_719 : _T_726;
  assign _T_728 = {_T_712,_T_727};
  assign _T_729 = _T_706[7:4];
  assign _T_730 = _T_706[3:0];
  assign _T_732 = _T_729 != 4'h0;
  assign _T_733 = _T_729[3];
  assign _T_735 = _T_729[2];
  assign _T_737 = _T_729[1];
  assign _T_738 = _T_735 ? 2'h2 : {{1'd0}, _T_737};
  assign _T_739 = _T_733 ? 2'h3 : _T_738;
  assign _T_740 = _T_730[3];
  assign _T_742 = _T_730[2];
  assign _T_744 = _T_730[1];
  assign _T_745 = _T_742 ? 2'h2 : {{1'd0}, _T_744};
  assign _T_746 = _T_740 ? 2'h3 : _T_745;
  assign _T_747 = _T_732 ? _T_739 : _T_746;
  assign _T_748 = {_T_732,_T_747};
  assign _T_749 = _T_708 ? _T_728 : _T_748;
  assign _T_750 = {_T_708,_T_749};
  assign _T_751 = _T_658 ? _T_704 : _T_750;
  assign _T_752 = {_T_658,_T_751};
  assign _T_753 = _T_556 ? _T_654 : _T_752;
  assign _T_754 = {_T_556,_T_753};
  assign _T_755 = _T_550[63:32];
  assign _T_756 = _T_550[31:0];
  assign _T_758 = _T_755 != 32'h0;
  assign _T_759 = _T_755[31:16];
  assign _T_760 = _T_755[15:0];
  assign _T_762 = _T_759 != 16'h0;
  assign _T_763 = _T_759[15:8];
  assign _T_764 = _T_759[7:0];
  assign _T_766 = _T_763 != 8'h0;
  assign _T_767 = _T_763[7:4];
  assign _T_768 = _T_763[3:0];
  assign _T_770 = _T_767 != 4'h0;
  assign _T_771 = _T_767[3];
  assign _T_773 = _T_767[2];
  assign _T_775 = _T_767[1];
  assign _T_776 = _T_773 ? 2'h2 : {{1'd0}, _T_775};
  assign _T_777 = _T_771 ? 2'h3 : _T_776;
  assign _T_778 = _T_768[3];
  assign _T_780 = _T_768[2];
  assign _T_782 = _T_768[1];
  assign _T_783 = _T_780 ? 2'h2 : {{1'd0}, _T_782};
  assign _T_784 = _T_778 ? 2'h3 : _T_783;
  assign _T_785 = _T_770 ? _T_777 : _T_784;
  assign _T_786 = {_T_770,_T_785};
  assign _T_787 = _T_764[7:4];
  assign _T_788 = _T_764[3:0];
  assign _T_790 = _T_787 != 4'h0;
  assign _T_791 = _T_787[3];
  assign _T_793 = _T_787[2];
  assign _T_795 = _T_787[1];
  assign _T_796 = _T_793 ? 2'h2 : {{1'd0}, _T_795};
  assign _T_797 = _T_791 ? 2'h3 : _T_796;
  assign _T_798 = _T_788[3];
  assign _T_800 = _T_788[2];
  assign _T_802 = _T_788[1];
  assign _T_803 = _T_800 ? 2'h2 : {{1'd0}, _T_802};
  assign _T_804 = _T_798 ? 2'h3 : _T_803;
  assign _T_805 = _T_790 ? _T_797 : _T_804;
  assign _T_806 = {_T_790,_T_805};
  assign _T_807 = _T_766 ? _T_786 : _T_806;
  assign _T_808 = {_T_766,_T_807};
  assign _T_809 = _T_760[15:8];
  assign _T_810 = _T_760[7:0];
  assign _T_812 = _T_809 != 8'h0;
  assign _T_813 = _T_809[7:4];
  assign _T_814 = _T_809[3:0];
  assign _T_816 = _T_813 != 4'h0;
  assign _T_817 = _T_813[3];
  assign _T_819 = _T_813[2];
  assign _T_821 = _T_813[1];
  assign _T_822 = _T_819 ? 2'h2 : {{1'd0}, _T_821};
  assign _T_823 = _T_817 ? 2'h3 : _T_822;
  assign _T_824 = _T_814[3];
  assign _T_826 = _T_814[2];
  assign _T_828 = _T_814[1];
  assign _T_829 = _T_826 ? 2'h2 : {{1'd0}, _T_828};
  assign _T_830 = _T_824 ? 2'h3 : _T_829;
  assign _T_831 = _T_816 ? _T_823 : _T_830;
  assign _T_832 = {_T_816,_T_831};
  assign _T_833 = _T_810[7:4];
  assign _T_834 = _T_810[3:0];
  assign _T_836 = _T_833 != 4'h0;
  assign _T_837 = _T_833[3];
  assign _T_839 = _T_833[2];
  assign _T_841 = _T_833[1];
  assign _T_842 = _T_839 ? 2'h2 : {{1'd0}, _T_841};
  assign _T_843 = _T_837 ? 2'h3 : _T_842;
  assign _T_844 = _T_834[3];
  assign _T_846 = _T_834[2];
  assign _T_848 = _T_834[1];
  assign _T_849 = _T_846 ? 2'h2 : {{1'd0}, _T_848};
  assign _T_850 = _T_844 ? 2'h3 : _T_849;
  assign _T_851 = _T_836 ? _T_843 : _T_850;
  assign _T_852 = {_T_836,_T_851};
  assign _T_853 = _T_812 ? _T_832 : _T_852;
  assign _T_854 = {_T_812,_T_853};
  assign _T_855 = _T_762 ? _T_808 : _T_854;
  assign _T_856 = {_T_762,_T_855};
  assign _T_857 = _T_756[31:16];
  assign _T_858 = _T_756[15:0];
  assign _T_860 = _T_857 != 16'h0;
  assign _T_861 = _T_857[15:8];
  assign _T_862 = _T_857[7:0];
  assign _T_864 = _T_861 != 8'h0;
  assign _T_865 = _T_861[7:4];
  assign _T_866 = _T_861[3:0];
  assign _T_868 = _T_865 != 4'h0;
  assign _T_869 = _T_865[3];
  assign _T_871 = _T_865[2];
  assign _T_873 = _T_865[1];
  assign _T_874 = _T_871 ? 2'h2 : {{1'd0}, _T_873};
  assign _T_875 = _T_869 ? 2'h3 : _T_874;
  assign _T_876 = _T_866[3];
  assign _T_878 = _T_866[2];
  assign _T_880 = _T_866[1];
  assign _T_881 = _T_878 ? 2'h2 : {{1'd0}, _T_880};
  assign _T_882 = _T_876 ? 2'h3 : _T_881;
  assign _T_883 = _T_868 ? _T_875 : _T_882;
  assign _T_884 = {_T_868,_T_883};
  assign _T_885 = _T_862[7:4];
  assign _T_886 = _T_862[3:0];
  assign _T_888 = _T_885 != 4'h0;
  assign _T_889 = _T_885[3];
  assign _T_891 = _T_885[2];
  assign _T_893 = _T_885[1];
  assign _T_894 = _T_891 ? 2'h2 : {{1'd0}, _T_893};
  assign _T_895 = _T_889 ? 2'h3 : _T_894;
  assign _T_896 = _T_886[3];
  assign _T_898 = _T_886[2];
  assign _T_900 = _T_886[1];
  assign _T_901 = _T_898 ? 2'h2 : {{1'd0}, _T_900};
  assign _T_902 = _T_896 ? 2'h3 : _T_901;
  assign _T_903 = _T_888 ? _T_895 : _T_902;
  assign _T_904 = {_T_888,_T_903};
  assign _T_905 = _T_864 ? _T_884 : _T_904;
  assign _T_906 = {_T_864,_T_905};
  assign _T_907 = _T_858[15:8];
  assign _T_908 = _T_858[7:0];
  assign _T_910 = _T_907 != 8'h0;
  assign _T_911 = _T_907[7:4];
  assign _T_912 = _T_907[3:0];
  assign _T_914 = _T_911 != 4'h0;
  assign _T_915 = _T_911[3];
  assign _T_917 = _T_911[2];
  assign _T_919 = _T_911[1];
  assign _T_920 = _T_917 ? 2'h2 : {{1'd0}, _T_919};
  assign _T_921 = _T_915 ? 2'h3 : _T_920;
  assign _T_922 = _T_912[3];
  assign _T_924 = _T_912[2];
  assign _T_926 = _T_912[1];
  assign _T_927 = _T_924 ? 2'h2 : {{1'd0}, _T_926};
  assign _T_928 = _T_922 ? 2'h3 : _T_927;
  assign _T_929 = _T_914 ? _T_921 : _T_928;
  assign _T_930 = {_T_914,_T_929};
  assign _T_931 = _T_908[7:4];
  assign _T_932 = _T_908[3:0];
  assign _T_934 = _T_931 != 4'h0;
  assign _T_935 = _T_931[3];
  assign _T_937 = _T_931[2];
  assign _T_939 = _T_931[1];
  assign _T_940 = _T_937 ? 2'h2 : {{1'd0}, _T_939};
  assign _T_941 = _T_935 ? 2'h3 : _T_940;
  assign _T_942 = _T_932[3];
  assign _T_944 = _T_932[2];
  assign _T_946 = _T_932[1];
  assign _T_947 = _T_944 ? 2'h2 : {{1'd0}, _T_946};
  assign _T_948 = _T_942 ? 2'h3 : _T_947;
  assign _T_949 = _T_934 ? _T_941 : _T_948;
  assign _T_950 = {_T_934,_T_949};
  assign _T_951 = _T_910 ? _T_930 : _T_950;
  assign _T_952 = {_T_910,_T_951};
  assign _T_953 = _T_860 ? _T_906 : _T_952;
  assign _T_954 = {_T_860,_T_953};
  assign _T_955 = _T_758 ? _T_856 : _T_954;
  assign _T_956 = {_T_758,_T_955};
  assign _T_957 = _T_552 ? _T_754 : _T_956;
  assign _T_958 = {_T_552,_T_957};
  assign _T_959 = _T_346 ? {{1'd0}, _T_548} : _T_958;
  assign _T_960 = {_T_346,_T_959};
  assign whichInterrupt = _T_960[4:0];
  assign _GEN_3 = {{27'd0}, whichInterrupt};
  assign _T_962 = 32'h80000000 + _GEN_3;
  assign interruptCause = _T_962[31:0];
  assign _T_964 = reg_debug == 1'h0;
  assign _T_965 = anyInterrupt & _T_964;
  assign _T_967 = io_singleStep == 1'h0;
  assign _T_968 = _T_965 & _T_967;
  assign _T_969 = _T_968 | reg_singleStepped;
  assign _T_971_mask = _T_982[31:0];
  assign _T_972 = reg_pmp_0_cfg_a[0];
  assign _T_973 = {reg_pmp_0_addr,_T_972};
  assign _T_977 = _T_973 + 31'h1;
  assign _T_978 = _T_977[30:0];
  assign _T_979 = ~ _T_978;
  assign _T_980 = _T_973 & _T_979;
  assign _T_982 = {_T_980,2'h3};
  assign _T_984_mask = _T_995[31:0];
  assign _T_985 = reg_pmp_1_cfg_a[0];
  assign _T_986 = {reg_pmp_1_addr,_T_985};
  assign _T_990 = _T_986 + 31'h1;
  assign _T_991 = _T_990[30:0];
  assign _T_992 = ~ _T_991;
  assign _T_993 = _T_986 & _T_992;
  assign _T_995 = {_T_993,2'h3};
  assign _T_997_mask = _T_1008[31:0];
  assign _T_998 = reg_pmp_2_cfg_a[0];
  assign _T_999 = {reg_pmp_2_addr,_T_998};
  assign _T_1003 = _T_999 + 31'h1;
  assign _T_1004 = _T_1003[30:0];
  assign _T_1005 = ~ _T_1004;
  assign _T_1006 = _T_999 & _T_1005;
  assign _T_1008 = {_T_1006,2'h3};
  assign _T_1010_mask = _T_1021[31:0];
  assign _T_1011 = reg_pmp_3_cfg_a[0];
  assign _T_1012 = {reg_pmp_3_addr,_T_1011};
  assign _T_1016 = _T_1012 + 31'h1;
  assign _T_1017 = _T_1016[30:0];
  assign _T_1018 = ~ _T_1017;
  assign _T_1019 = _T_1012 & _T_1018;
  assign _T_1021 = {_T_1019,2'h3};
  assign _T_1023_mask = _T_1034[31:0];
  assign _T_1024 = reg_pmp_4_cfg_a[0];
  assign _T_1025 = {reg_pmp_4_addr,_T_1024};
  assign _T_1029 = _T_1025 + 31'h1;
  assign _T_1030 = _T_1029[30:0];
  assign _T_1031 = ~ _T_1030;
  assign _T_1032 = _T_1025 & _T_1031;
  assign _T_1034 = {_T_1032,2'h3};
  assign _T_1036_mask = _T_1047[31:0];
  assign _T_1037 = reg_pmp_5_cfg_a[0];
  assign _T_1038 = {reg_pmp_5_addr,_T_1037};
  assign _T_1042 = _T_1038 + 31'h1;
  assign _T_1043 = _T_1042[30:0];
  assign _T_1044 = ~ _T_1043;
  assign _T_1045 = _T_1038 & _T_1044;
  assign _T_1047 = {_T_1045,2'h3};
  assign _T_1049_mask = _T_1060[31:0];
  assign _T_1050 = reg_pmp_6_cfg_a[0];
  assign _T_1051 = {reg_pmp_6_addr,_T_1050};
  assign _T_1055 = _T_1051 + 31'h1;
  assign _T_1056 = _T_1055[30:0];
  assign _T_1057 = ~ _T_1056;
  assign _T_1058 = _T_1051 & _T_1057;
  assign _T_1060 = {_T_1058,2'h3};
  assign _T_1062_mask = _T_1073[31:0];
  assign _T_1063 = reg_pmp_7_cfg_a[0];
  assign _T_1064 = {reg_pmp_7_addr,_T_1063};
  assign _T_1068 = _T_1064 + 31'h1;
  assign _T_1069 = _T_1068[30:0];
  assign _T_1070 = ~ _T_1069;
  assign _T_1071 = _T_1064 & _T_1070;
  assign _T_1073 = {_T_1071,2'h3};
  assign _T_1076 = {io_status_hie,io_status_sie};
  assign _T_1077 = {_T_1076,io_status_uie};
  assign _T_1078 = {io_status_upie,io_status_mie};
  assign _T_1079 = {io_status_hpie,io_status_spie};
  assign _T_1080 = {_T_1079,_T_1078};
  assign _T_1081 = {_T_1080,_T_1077};
  assign _T_1082 = {io_status_hpp,io_status_spp};
  assign _T_1083 = {_T_1082,io_status_mpie};
  assign _T_1084 = {io_status_fs,io_status_mpp};
  assign _T_1085 = {io_status_mprv,io_status_xs};
  assign _T_1086 = {_T_1085,_T_1084};
  assign _T_1087 = {_T_1086,_T_1083};
  assign _T_1088 = {_T_1087,_T_1081};
  assign _T_1089 = {io_status_tvm,io_status_mxr};
  assign _T_1090 = {_T_1089,io_status_sum};
  assign _T_1091 = {io_status_tsr,io_status_tw};
  assign _T_1092 = {io_status_sd_rv32,io_status_zero1};
  assign _T_1093 = {_T_1092,_T_1091};
  assign _T_1094 = {_T_1093,_T_1090};
  assign _T_1095 = {io_status_sxl,io_status_uxl};
  assign _T_1096 = {io_status_sd,io_status_zero2};
  assign _T_1097 = {_T_1096,_T_1095};
  assign _T_1098 = {io_status_dprv,io_status_prv};
  assign _T_1099 = {io_status_debug,io_status_isa};
  assign _T_1100 = {_T_1099,_T_1098};
  assign _T_1101 = {_T_1100,_T_1097};
  assign _T_1102 = {_T_1101,_T_1094};
  assign _T_1103 = {_T_1102,_T_1088};
  assign read_mstatus = _T_1103[31:0];
  assign _GEN_37 = reg_tselect ? reg_bp_1_control_ttype : reg_bp_0_control_ttype;
  assign _GEN_38 = reg_tselect ? reg_bp_1_control_dmode : reg_bp_0_control_dmode;
  assign _GEN_39 = reg_tselect ? reg_bp_1_control_maskmax : reg_bp_0_control_maskmax;
  assign _GEN_40 = reg_tselect ? reg_bp_1_control_reserved : reg_bp_0_control_reserved;
  assign _GEN_41 = reg_tselect ? reg_bp_1_control_action : reg_bp_0_control_action;
  assign _GEN_42 = reg_tselect ? reg_bp_1_control_chain : reg_bp_0_control_chain;
  assign _GEN_43 = reg_tselect ? reg_bp_1_control_zero : reg_bp_0_control_zero;
  assign _GEN_44 = reg_tselect ? reg_bp_1_control_tmatch : reg_bp_0_control_tmatch;
  assign _GEN_45 = reg_tselect ? reg_bp_1_control_m : reg_bp_0_control_m;
  assign _GEN_46 = reg_tselect ? reg_bp_1_control_h : reg_bp_0_control_h;
  assign _GEN_47 = reg_tselect ? reg_bp_1_control_s : reg_bp_0_control_s;
  assign _GEN_48 = reg_tselect ? reg_bp_1_control_u : reg_bp_0_control_u;
  assign _GEN_49 = reg_tselect ? reg_bp_1_control_x : reg_bp_0_control_x;
  assign _GEN_50 = reg_tselect ? reg_bp_1_control_w : reg_bp_0_control_w;
  assign _GEN_51 = reg_tselect ? reg_bp_1_control_r : reg_bp_0_control_r;
  assign _GEN_52 = reg_tselect ? reg_bp_1_address : reg_bp_0_address;
  assign _T_1105 = {_GEN_49,_GEN_50};
  assign _T_1106 = {_T_1105,_GEN_51};
  assign _T_1107 = {_GEN_47,_GEN_48};
  assign _T_1108 = {_GEN_45,_GEN_46};
  assign _T_1109 = {_T_1108,_T_1107};
  assign _T_1110 = {_T_1109,_T_1106};
  assign _T_1111 = {_GEN_43,_GEN_44};
  assign _T_1112 = {_GEN_41,_GEN_42};
  assign _T_1113 = {_T_1112,_T_1111};
  assign _T_1114 = {_GEN_39,_GEN_40};
  assign _T_1115 = {_GEN_37,_GEN_38};
  assign _T_1116 = {_T_1115,_T_1114};
  assign _T_1117 = {_T_1116,_T_1113};
  assign _T_1118 = {_T_1117,_T_1110};
  assign _T_1123 = {reg_dcsr_zero1,reg_dcsr_step};
  assign _T_1124 = {_T_1123,reg_dcsr_prv};
  assign _T_1125 = {reg_dcsr_stoptime,reg_dcsr_cause};
  assign _T_1126 = {reg_dcsr_zero2,reg_dcsr_stopcycle};
  assign _T_1127 = {_T_1126,_T_1125};
  assign _T_1128 = {_T_1127,_T_1124};
  assign _T_1129 = {reg_dcsr_ebreakh,reg_dcsr_ebreaks};
  assign _T_1130 = {_T_1129,reg_dcsr_ebreaku};
  assign _T_1131 = {reg_dcsr_zero3,reg_dcsr_ebreakm};
  assign _T_1132 = {reg_dcsr_xdebugver,reg_dcsr_zero4};
  assign _T_1133 = {_T_1132,_T_1131};
  assign _T_1134 = {_T_1133,_T_1130};
  assign _T_1135 = {_T_1134,_T_1128};
  assign _T_1139 = _T_270[63:32];
  assign _T_1140 = _T_257[63:32];
  assign _T_1156 = {reg_pmp_0_cfg_x,reg_pmp_0_cfg_w};
  assign _T_1157 = {_T_1156,reg_pmp_0_cfg_r};
  assign _T_1158 = {reg_pmp_0_cfg_l,reg_pmp_0_cfg_res};
  assign _T_1159 = {_T_1158,reg_pmp_0_cfg_a};
  assign _T_1160 = {_T_1159,_T_1157};
  assign _T_1161 = {reg_pmp_1_cfg_x,reg_pmp_1_cfg_w};
  assign _T_1162 = {_T_1161,reg_pmp_1_cfg_r};
  assign _T_1163 = {reg_pmp_1_cfg_l,reg_pmp_1_cfg_res};
  assign _T_1164 = {_T_1163,reg_pmp_1_cfg_a};
  assign _T_1165 = {_T_1164,_T_1162};
  assign _T_1166 = {reg_pmp_2_cfg_x,reg_pmp_2_cfg_w};
  assign _T_1167 = {_T_1166,reg_pmp_2_cfg_r};
  assign _T_1168 = {reg_pmp_2_cfg_l,reg_pmp_2_cfg_res};
  assign _T_1169 = {_T_1168,reg_pmp_2_cfg_a};
  assign _T_1170 = {_T_1169,_T_1167};
  assign _T_1171 = {reg_pmp_3_cfg_x,reg_pmp_3_cfg_w};
  assign _T_1172 = {_T_1171,reg_pmp_3_cfg_r};
  assign _T_1173 = {reg_pmp_3_cfg_l,reg_pmp_3_cfg_res};
  assign _T_1174 = {_T_1173,reg_pmp_3_cfg_a};
  assign _T_1175 = {_T_1174,_T_1172};
  assign _T_1176 = {_T_1165,_T_1160};
  assign _T_1177 = {_T_1175,_T_1170};
  assign _T_1178 = {_T_1177,_T_1176};
  assign _T_1179 = {reg_pmp_4_cfg_x,reg_pmp_4_cfg_w};
  assign _T_1180 = {_T_1179,reg_pmp_4_cfg_r};
  assign _T_1181 = {reg_pmp_4_cfg_l,reg_pmp_4_cfg_res};
  assign _T_1182 = {_T_1181,reg_pmp_4_cfg_a};
  assign _T_1183 = {_T_1182,_T_1180};
  assign _T_1184 = {reg_pmp_5_cfg_x,reg_pmp_5_cfg_w};
  assign _T_1185 = {_T_1184,reg_pmp_5_cfg_r};
  assign _T_1186 = {reg_pmp_5_cfg_l,reg_pmp_5_cfg_res};
  assign _T_1187 = {_T_1186,reg_pmp_5_cfg_a};
  assign _T_1188 = {_T_1187,_T_1185};
  assign _T_1189 = {reg_pmp_6_cfg_x,reg_pmp_6_cfg_w};
  assign _T_1190 = {_T_1189,reg_pmp_6_cfg_r};
  assign _T_1191 = {reg_pmp_6_cfg_l,reg_pmp_6_cfg_res};
  assign _T_1192 = {_T_1191,reg_pmp_6_cfg_a};
  assign _T_1193 = {_T_1192,_T_1190};
  assign _T_1194 = {reg_pmp_7_cfg_x,reg_pmp_7_cfg_w};
  assign _T_1195 = {_T_1194,reg_pmp_7_cfg_r};
  assign _T_1196 = {reg_pmp_7_cfg_l,reg_pmp_7_cfg_res};
  assign _T_1197 = {_T_1196,reg_pmp_7_cfg_a};
  assign _T_1198 = {_T_1197,_T_1195};
  assign _T_1199 = {_T_1188,_T_1183};
  assign _T_1200 = {_T_1198,_T_1193};
  assign _T_1201 = {_T_1200,_T_1199};
  assign _T_1249 = io_rw_addr == 12'h7a0;
  assign _T_1251 = io_rw_addr == 12'h7a1;
  assign _T_1253 = io_rw_addr == 12'h7a2;
  assign _T_1261 = io_rw_addr == 12'hb00;
  assign _T_1263 = io_rw_addr == 12'hb02;
  assign _T_1265 = io_rw_addr == 12'h301;
  assign _T_1267 = io_rw_addr == 12'h300;
  assign _T_1269 = io_rw_addr == 12'h305;
  assign _T_1271 = io_rw_addr == 12'h344;
  assign _T_1273 = io_rw_addr == 12'h304;
  assign _T_1275 = io_rw_addr == 12'h340;
  assign _T_1277 = io_rw_addr == 12'h341;
  assign _T_1279 = io_rw_addr == 12'h343;
  assign _T_1281 = io_rw_addr == 12'h342;
  assign _T_1283 = io_rw_addr == 12'hf14;
  assign _T_1285 = io_rw_addr == 12'h7b0;
  assign _T_1287 = io_rw_addr == 12'h7b1;
  assign _T_1289 = io_rw_addr == 12'h7b2;
  assign _T_1465 = io_rw_addr == 12'hb80;
  assign _T_1467 = io_rw_addr == 12'hb82;
  assign _T_1469 = io_rw_addr == 12'h3a0;
  assign _T_1471 = io_rw_addr == 12'h3a1;
  assign _T_1477 = io_rw_addr == 12'h3b0;
  assign _T_1479 = io_rw_addr == 12'h3b1;
  assign _T_1481 = io_rw_addr == 12'h3b2;
  assign _T_1483 = io_rw_addr == 12'h3b3;
  assign _T_1485 = io_rw_addr == 12'h3b4;
  assign _T_1487 = io_rw_addr == 12'h3b5;
  assign _T_1489 = io_rw_addr == 12'h3b6;
  assign _T_1491 = io_rw_addr == 12'h3b7;
  assign _T_1510 = io_rw_cmd == 3'h2;
  assign _T_1511 = io_rw_cmd == 3'h3;
  assign _T_1512 = _T_1510 | _T_1511;
  assign _T_1514 = _T_1512 ? io_rw_rdata : 32'h0;
  assign _T_1515 = _T_1514 | io_rw_wdata;
  assign _T_1519 = _T_1511 ? io_rw_wdata : 32'h0;
  assign _T_1520 = ~ _T_1519;
  assign wdata = _T_1515 & _T_1520;
  assign system_insn = io_rw_cmd == 3'h4;
  assign _T_1523 = io_rw_addr[2:0];
  assign opcode = 8'h1 << _T_1523;
  assign _T_1524 = opcode[0];
  assign insn_call = system_insn & _T_1524;
  assign _T_1525 = opcode[1];
  assign insn_break = system_insn & _T_1525;
  assign _T_1526 = opcode[2];
  assign insn_ret = system_insn & _T_1526;
  assign _T_1527 = opcode[5];
  assign insn_wfi = system_insn & _T_1527;
  assign _T_1558 = io_decode_csr[9:8];
  assign _T_1559 = reg_mstatus_prv < _T_1558;
  assign _T_1561 = io_decode_csr == 12'h7a0;
  assign _T_1563 = io_decode_csr == 12'h7a1;
  assign _T_1565 = io_decode_csr == 12'h7a2;
  assign _T_1567 = io_decode_csr == 12'hf13;
  assign _T_1569 = io_decode_csr == 12'hf12;
  assign _T_1571 = io_decode_csr == 12'hf11;
  assign _T_1573 = io_decode_csr == 12'hb00;
  assign _T_1575 = io_decode_csr == 12'hb02;
  assign _T_1577 = io_decode_csr == 12'h301;
  assign _T_1579 = io_decode_csr == 12'h300;
  assign _T_1581 = io_decode_csr == 12'h305;
  assign _T_1583 = io_decode_csr == 12'h344;
  assign _T_1585 = io_decode_csr == 12'h304;
  assign _T_1587 = io_decode_csr == 12'h340;
  assign _T_1589 = io_decode_csr == 12'h341;
  assign _T_1591 = io_decode_csr == 12'h343;
  assign _T_1593 = io_decode_csr == 12'h342;
  assign _T_1595 = io_decode_csr == 12'hf14;
  assign _T_1597 = io_decode_csr == 12'h7b0;
  assign _T_1599 = io_decode_csr == 12'h7b1;
  assign _T_1601 = io_decode_csr == 12'h7b2;
  assign _T_1603 = io_decode_csr == 12'h323;
  assign _T_1605 = io_decode_csr == 12'hb03;
  assign _T_1607 = io_decode_csr == 12'hb83;
  assign _T_1609 = io_decode_csr == 12'h324;
  assign _T_1611 = io_decode_csr == 12'hb04;
  assign _T_1613 = io_decode_csr == 12'hb84;
  assign _T_1615 = io_decode_csr == 12'h325;
  assign _T_1617 = io_decode_csr == 12'hb05;
  assign _T_1619 = io_decode_csr == 12'hb85;
  assign _T_1621 = io_decode_csr == 12'h326;
  assign _T_1623 = io_decode_csr == 12'hb06;
  assign _T_1625 = io_decode_csr == 12'hb86;
  assign _T_1627 = io_decode_csr == 12'h327;
  assign _T_1629 = io_decode_csr == 12'hb07;
  assign _T_1631 = io_decode_csr == 12'hb87;
  assign _T_1633 = io_decode_csr == 12'h328;
  assign _T_1635 = io_decode_csr == 12'hb08;
  assign _T_1637 = io_decode_csr == 12'hb88;
  assign _T_1639 = io_decode_csr == 12'h329;
  assign _T_1641 = io_decode_csr == 12'hb09;
  assign _T_1643 = io_decode_csr == 12'hb89;
  assign _T_1645 = io_decode_csr == 12'h32a;
  assign _T_1647 = io_decode_csr == 12'hb0a;
  assign _T_1649 = io_decode_csr == 12'hb8a;
  assign _T_1651 = io_decode_csr == 12'h32b;
  assign _T_1653 = io_decode_csr == 12'hb0b;
  assign _T_1655 = io_decode_csr == 12'hb8b;
  assign _T_1657 = io_decode_csr == 12'h32c;
  assign _T_1659 = io_decode_csr == 12'hb0c;
  assign _T_1661 = io_decode_csr == 12'hb8c;
  assign _T_1663 = io_decode_csr == 12'h32d;
  assign _T_1665 = io_decode_csr == 12'hb0d;
  assign _T_1667 = io_decode_csr == 12'hb8d;
  assign _T_1669 = io_decode_csr == 12'h32e;
  assign _T_1671 = io_decode_csr == 12'hb0e;
  assign _T_1673 = io_decode_csr == 12'hb8e;
  assign _T_1675 = io_decode_csr == 12'h32f;
  assign _T_1677 = io_decode_csr == 12'hb0f;
  assign _T_1679 = io_decode_csr == 12'hb8f;
  assign _T_1681 = io_decode_csr == 12'h330;
  assign _T_1683 = io_decode_csr == 12'hb10;
  assign _T_1685 = io_decode_csr == 12'hb90;
  assign _T_1687 = io_decode_csr == 12'h331;
  assign _T_1689 = io_decode_csr == 12'hb11;
  assign _T_1691 = io_decode_csr == 12'hb91;
  assign _T_1693 = io_decode_csr == 12'h332;
  assign _T_1695 = io_decode_csr == 12'hb12;
  assign _T_1697 = io_decode_csr == 12'hb92;
  assign _T_1699 = io_decode_csr == 12'h333;
  assign _T_1701 = io_decode_csr == 12'hb13;
  assign _T_1703 = io_decode_csr == 12'hb93;
  assign _T_1705 = io_decode_csr == 12'h334;
  assign _T_1707 = io_decode_csr == 12'hb14;
  assign _T_1709 = io_decode_csr == 12'hb94;
  assign _T_1711 = io_decode_csr == 12'h335;
  assign _T_1713 = io_decode_csr == 12'hb15;
  assign _T_1715 = io_decode_csr == 12'hb95;
  assign _T_1717 = io_decode_csr == 12'h336;
  assign _T_1719 = io_decode_csr == 12'hb16;
  assign _T_1721 = io_decode_csr == 12'hb96;
  assign _T_1723 = io_decode_csr == 12'h337;
  assign _T_1725 = io_decode_csr == 12'hb17;
  assign _T_1727 = io_decode_csr == 12'hb97;
  assign _T_1729 = io_decode_csr == 12'h338;
  assign _T_1731 = io_decode_csr == 12'hb18;
  assign _T_1733 = io_decode_csr == 12'hb98;
  assign _T_1735 = io_decode_csr == 12'h339;
  assign _T_1737 = io_decode_csr == 12'hb19;
  assign _T_1739 = io_decode_csr == 12'hb99;
  assign _T_1741 = io_decode_csr == 12'h33a;
  assign _T_1743 = io_decode_csr == 12'hb1a;
  assign _T_1745 = io_decode_csr == 12'hb9a;
  assign _T_1747 = io_decode_csr == 12'h33b;
  assign _T_1749 = io_decode_csr == 12'hb1b;
  assign _T_1751 = io_decode_csr == 12'hb9b;
  assign _T_1753 = io_decode_csr == 12'h33c;
  assign _T_1755 = io_decode_csr == 12'hb1c;
  assign _T_1757 = io_decode_csr == 12'hb9c;
  assign _T_1759 = io_decode_csr == 12'h33d;
  assign _T_1761 = io_decode_csr == 12'hb1d;
  assign _T_1763 = io_decode_csr == 12'hb9d;
  assign _T_1765 = io_decode_csr == 12'h33e;
  assign _T_1767 = io_decode_csr == 12'hb1e;
  assign _T_1769 = io_decode_csr == 12'hb9e;
  assign _T_1771 = io_decode_csr == 12'h33f;
  assign _T_1773 = io_decode_csr == 12'hb1f;
  assign _T_1775 = io_decode_csr == 12'hb9f;
  assign _T_1777 = io_decode_csr == 12'hb80;
  assign _T_1779 = io_decode_csr == 12'hb82;
  assign _T_1781 = io_decode_csr == 12'h3a0;
  assign _T_1783 = io_decode_csr == 12'h3a1;
  assign _T_1785 = io_decode_csr == 12'h3a2;
  assign _T_1787 = io_decode_csr == 12'h3a3;
  assign _T_1789 = io_decode_csr == 12'h3b0;
  assign _T_1791 = io_decode_csr == 12'h3b1;
  assign _T_1793 = io_decode_csr == 12'h3b2;
  assign _T_1795 = io_decode_csr == 12'h3b3;
  assign _T_1797 = io_decode_csr == 12'h3b4;
  assign _T_1799 = io_decode_csr == 12'h3b5;
  assign _T_1801 = io_decode_csr == 12'h3b6;
  assign _T_1803 = io_decode_csr == 12'h3b7;
  assign _T_1805 = io_decode_csr == 12'h3b8;
  assign _T_1807 = io_decode_csr == 12'h3b9;
  assign _T_1809 = io_decode_csr == 12'h3ba;
  assign _T_1811 = io_decode_csr == 12'h3bb;
  assign _T_1813 = io_decode_csr == 12'h3bc;
  assign _T_1815 = io_decode_csr == 12'h3bd;
  assign _T_1817 = io_decode_csr == 12'h3be;
  assign _T_1819 = io_decode_csr == 12'h3bf;
  assign _T_1820 = _T_1561 | _T_1563;
  assign _T_1821 = _T_1820 | _T_1565;
  assign _T_1822 = _T_1821 | _T_1567;
  assign _T_1823 = _T_1822 | _T_1569;
  assign _T_1824 = _T_1823 | _T_1571;
  assign _T_1825 = _T_1824 | _T_1573;
  assign _T_1826 = _T_1825 | _T_1575;
  assign _T_1827 = _T_1826 | _T_1577;
  assign _T_1828 = _T_1827 | _T_1579;
  assign _T_1829 = _T_1828 | _T_1581;
  assign _T_1830 = _T_1829 | _T_1583;
  assign _T_1831 = _T_1830 | _T_1585;
  assign _T_1832 = _T_1831 | _T_1587;
  assign _T_1833 = _T_1832 | _T_1589;
  assign _T_1834 = _T_1833 | _T_1591;
  assign _T_1835 = _T_1834 | _T_1593;
  assign _T_1836 = _T_1835 | _T_1595;
  assign _T_1837 = _T_1836 | _T_1597;
  assign _T_1838 = _T_1837 | _T_1599;
  assign _T_1839 = _T_1838 | _T_1601;
  assign _T_1840 = _T_1839 | _T_1603;
  assign _T_1841 = _T_1840 | _T_1605;
  assign _T_1842 = _T_1841 | _T_1607;
  assign _T_1843 = _T_1842 | _T_1609;
  assign _T_1844 = _T_1843 | _T_1611;
  assign _T_1845 = _T_1844 | _T_1613;
  assign _T_1846 = _T_1845 | _T_1615;
  assign _T_1847 = _T_1846 | _T_1617;
  assign _T_1848 = _T_1847 | _T_1619;
  assign _T_1849 = _T_1848 | _T_1621;
  assign _T_1850 = _T_1849 | _T_1623;
  assign _T_1851 = _T_1850 | _T_1625;
  assign _T_1852 = _T_1851 | _T_1627;
  assign _T_1853 = _T_1852 | _T_1629;
  assign _T_1854 = _T_1853 | _T_1631;
  assign _T_1855 = _T_1854 | _T_1633;
  assign _T_1856 = _T_1855 | _T_1635;
  assign _T_1857 = _T_1856 | _T_1637;
  assign _T_1858 = _T_1857 | _T_1639;
  assign _T_1859 = _T_1858 | _T_1641;
  assign _T_1860 = _T_1859 | _T_1643;
  assign _T_1861 = _T_1860 | _T_1645;
  assign _T_1862 = _T_1861 | _T_1647;
  assign _T_1863 = _T_1862 | _T_1649;
  assign _T_1864 = _T_1863 | _T_1651;
  assign _T_1865 = _T_1864 | _T_1653;
  assign _T_1866 = _T_1865 | _T_1655;
  assign _T_1867 = _T_1866 | _T_1657;
  assign _T_1868 = _T_1867 | _T_1659;
  assign _T_1869 = _T_1868 | _T_1661;
  assign _T_1870 = _T_1869 | _T_1663;
  assign _T_1871 = _T_1870 | _T_1665;
  assign _T_1872 = _T_1871 | _T_1667;
  assign _T_1873 = _T_1872 | _T_1669;
  assign _T_1874 = _T_1873 | _T_1671;
  assign _T_1875 = _T_1874 | _T_1673;
  assign _T_1876 = _T_1875 | _T_1675;
  assign _T_1877 = _T_1876 | _T_1677;
  assign _T_1878 = _T_1877 | _T_1679;
  assign _T_1879 = _T_1878 | _T_1681;
  assign _T_1880 = _T_1879 | _T_1683;
  assign _T_1881 = _T_1880 | _T_1685;
  assign _T_1882 = _T_1881 | _T_1687;
  assign _T_1883 = _T_1882 | _T_1689;
  assign _T_1884 = _T_1883 | _T_1691;
  assign _T_1885 = _T_1884 | _T_1693;
  assign _T_1886 = _T_1885 | _T_1695;
  assign _T_1887 = _T_1886 | _T_1697;
  assign _T_1888 = _T_1887 | _T_1699;
  assign _T_1889 = _T_1888 | _T_1701;
  assign _T_1890 = _T_1889 | _T_1703;
  assign _T_1891 = _T_1890 | _T_1705;
  assign _T_1892 = _T_1891 | _T_1707;
  assign _T_1893 = _T_1892 | _T_1709;
  assign _T_1894 = _T_1893 | _T_1711;
  assign _T_1895 = _T_1894 | _T_1713;
  assign _T_1896 = _T_1895 | _T_1715;
  assign _T_1897 = _T_1896 | _T_1717;
  assign _T_1898 = _T_1897 | _T_1719;
  assign _T_1899 = _T_1898 | _T_1721;
  assign _T_1900 = _T_1899 | _T_1723;
  assign _T_1901 = _T_1900 | _T_1725;
  assign _T_1902 = _T_1901 | _T_1727;
  assign _T_1903 = _T_1902 | _T_1729;
  assign _T_1904 = _T_1903 | _T_1731;
  assign _T_1905 = _T_1904 | _T_1733;
  assign _T_1906 = _T_1905 | _T_1735;
  assign _T_1907 = _T_1906 | _T_1737;
  assign _T_1908 = _T_1907 | _T_1739;
  assign _T_1909 = _T_1908 | _T_1741;
  assign _T_1910 = _T_1909 | _T_1743;
  assign _T_1911 = _T_1910 | _T_1745;
  assign _T_1912 = _T_1911 | _T_1747;
  assign _T_1913 = _T_1912 | _T_1749;
  assign _T_1914 = _T_1913 | _T_1751;
  assign _T_1915 = _T_1914 | _T_1753;
  assign _T_1916 = _T_1915 | _T_1755;
  assign _T_1917 = _T_1916 | _T_1757;
  assign _T_1918 = _T_1917 | _T_1759;
  assign _T_1919 = _T_1918 | _T_1761;
  assign _T_1920 = _T_1919 | _T_1763;
  assign _T_1921 = _T_1920 | _T_1765;
  assign _T_1922 = _T_1921 | _T_1767;
  assign _T_1923 = _T_1922 | _T_1769;
  assign _T_1924 = _T_1923 | _T_1771;
  assign _T_1925 = _T_1924 | _T_1773;
  assign _T_1926 = _T_1925 | _T_1775;
  assign _T_1927 = _T_1926 | _T_1777;
  assign _T_1928 = _T_1927 | _T_1779;
  assign _T_1929 = _T_1928 | _T_1781;
  assign _T_1930 = _T_1929 | _T_1783;
  assign _T_1931 = _T_1930 | _T_1785;
  assign _T_1932 = _T_1931 | _T_1787;
  assign _T_1933 = _T_1932 | _T_1789;
  assign _T_1934 = _T_1933 | _T_1791;
  assign _T_1935 = _T_1934 | _T_1793;
  assign _T_1936 = _T_1935 | _T_1795;
  assign _T_1937 = _T_1936 | _T_1797;
  assign _T_1938 = _T_1937 | _T_1799;
  assign _T_1939 = _T_1938 | _T_1801;
  assign _T_1940 = _T_1939 | _T_1803;
  assign _T_1941 = _T_1940 | _T_1805;
  assign _T_1942 = _T_1941 | _T_1807;
  assign _T_1943 = _T_1942 | _T_1809;
  assign _T_1944 = _T_1943 | _T_1811;
  assign _T_1945 = _T_1944 | _T_1813;
  assign _T_1946 = _T_1945 | _T_1815;
  assign _T_1947 = _T_1946 | _T_1817;
  assign _T_1948 = _T_1947 | _T_1819;
  assign _T_1950 = _T_1948 == 1'h0;
  assign _T_1951 = _T_1559 | _T_1950;
  assign _T_1960 = io_decode_csr >= 12'hc00;
  assign _T_1961 = io_decode_csr < 12'hc20;
  assign _T_1962 = _T_1960 & _T_1961;
  assign _T_1965 = io_decode_csr >= 12'hc80;
  assign _T_1966 = io_decode_csr < 12'hca0;
  assign _T_1967 = _T_1965 & _T_1966;
  assign _T_1968 = _T_1962 | _T_1967;
  assign _T_1971 = _T_1968 & _T_298;
  assign _T_1973 = hpm_mask >> io_decode_csr;
  assign _T_1974 = _T_1973[0];
  assign _T_1975 = _T_1971 & _T_1974;
  assign _T_1976 = _T_1951 | _T_1975;
  assign _T_1984 = _T_1597 | _T_1599;
  assign _T_1985 = _T_1984 | _T_1601;
  assign _T_1989 = _T_1985 & _T_964;
  assign _T_1990 = _T_1976 | _T_1989;
  assign _T_2003 = io_decode_csr[11:10];
  assign _T_2004 = ~ _T_2003;
  assign _T_2006 = _T_2004 == 2'h0;
  assign _T_2008 = io_decode_csr >= 12'h340;
  assign _T_2010 = io_decode_csr <= 12'h343;
  assign _T_2011 = _T_2008 & _T_2010;
  assign _T_2013 = io_decode_csr >= 12'h140;
  assign _T_2015 = io_decode_csr <= 12'h143;
  assign _T_2016 = _T_2013 & _T_2015;
  assign _T_2017 = _T_2011 | _T_2016;
  assign _T_2019 = _T_2017 == 1'h0;
  assign _GEN_4 = {{2'd0}, reg_mstatus_prv};
  assign _T_2046 = _GEN_4 + 4'h8;
  assign _T_2047 = _T_2046[3:0];
  assign _T_2049 = insn_break ? 32'h3 : io_cause;
  assign cause = insn_call ? {{28'd0}, _T_2047} : _T_2049;
  assign cause_lsbs = cause[4:0];
  assign _T_2050 = cause[31];
  assign _T_2052 = cause_lsbs == 5'he;
  assign causeIsDebugInt = _T_2050 & _T_2052;
  assign _T_2055 = _T_2050 == 1'h0;
  assign causeIsDebugTrigger = _T_2055 & _T_2052;
  assign _T_2061 = _T_2055 & insn_break;
  assign _T_2062 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign _T_2063 = {reg_dcsr_ebreakm,reg_dcsr_ebreakh};
  assign _T_2064 = {_T_2063,_T_2062};
  assign _T_2065 = _T_2064 >> reg_mstatus_prv;
  assign _T_2066 = _T_2065[0];
  assign causeIsDebugBreak = _T_2061 & _T_2066;
  assign _T_2068 = reg_singleStepped | causeIsDebugInt;
  assign _T_2069 = _T_2068 | causeIsDebugTrigger;
  assign _T_2070 = _T_2069 | causeIsDebugBreak;
  assign _T_2071 = _T_2070 | reg_debug;
  assign _T_2074 = insn_break ? 12'h800 : 12'h808;
  assign debugTVec = reg_debug ? _T_2074 : 12'h800;
  assign _T_2090 = cause[3:0];
  assign _GEN_5 = {{2'd0}, _T_2090};
  assign _T_2091 = _GEN_5 << 2;
  assign _T_2092 = reg_mtvec[31:6];
  assign _T_2093 = {_T_2092,_T_2091};
  assign _T_2094 = reg_mtvec[0];
  assign _T_2096 = _T_2094 & _T_2050;
  assign notDebugTVec = _T_2096 ? _T_2093 : reg_mtvec;
  assign tvec = _T_2071 ? {{20'd0}, debugTVec} : notDebugTVec;
  assign _T_2097 = insn_call | insn_break;
  assign _T_2098 = _T_2097 | insn_ret;
  assign _T_2101 = reg_dcsr_step & _T_964;
  assign _T_2102 = ~ io_status_fs;
  assign _T_2104 = _T_2102 == 2'h0;
  assign _T_2105 = ~ io_status_xs;
  assign _T_2107 = _T_2105 == 2'h0;
  assign _T_2108 = _T_2104 | _T_2107;
  assign _T_2113 = reg_mstatus_mprv & _T_964;
  assign _T_2114 = _T_2113 ? reg_mstatus_mpp : reg_mstatus_prv;
  assign exception = _T_2097 | io_exception;
  assign _T_2118 = insn_ret + insn_call;
  assign _T_2119 = insn_break + io_exception;
  assign _T_2120 = _T_2118 + _T_2119;
  assign _T_2122 = _T_2120 <= 3'h1;
  assign _T_2123 = _T_2122 | reset;
  assign _T_2125 = _T_2123 == 1'h0;
  assign _T_2128 = insn_wfi & _T_967;
  assign _T_2131 = _T_2128 & _T_964;
  assign _GEN_53 = _T_2131 ? 1'h1 : reg_wfi;
  assign _T_2134 = pending_interrupts != 32'h0;
  assign _T_2135 = _T_2134 | exception;
  assign _T_2136 = _T_2135 | reg_debugint;
  assign _GEN_54 = _T_2136 ? 1'h0 : _GEN_53;
  assign _T_2139 = reg_wfi == 1'h0;
  assign _T_2141 = io_retire == 1'h0;
  assign _T_2142 = _T_2139 | _T_2141;
  assign _T_2143 = _T_2142 | reset;
  assign _T_2145 = _T_2143 == 1'h0;
  assign _T_2147 = io_retire | exception;
  assign _GEN_55 = _T_2147 ? 1'h1 : reg_singleStepped;
  assign _GEN_56 = _T_967 ? 1'h0 : _GEN_55;
  assign _T_2161 = reg_singleStepped == 1'h0;
  assign _T_2164 = _T_2161 | _T_2141;
  assign _T_2165 = _T_2164 | reset;
  assign _T_2167 = _T_2165 == 1'h0;
  assign _T_2168 = ~ io_pc;
  assign _T_2170 = _T_2168 | 32'h1;
  assign _T_2171 = ~ _T_2170;
  assign _T_2183 = cause == 32'h2;
  assign _T_2184 = cause == 32'h3;
  assign _T_2185 = cause == 32'h4;
  assign _T_2186 = cause == 32'h6;
  assign _T_2187 = cause == 32'h0;
  assign _T_2188 = cause == 32'h5;
  assign _T_2189 = cause == 32'h7;
  assign _T_2190 = cause == 32'h1;
  assign _T_2191 = cause == 32'hd;
  assign _T_2192 = cause == 32'hf;
  assign _T_2193 = cause == 32'hc;
  assign _T_2194 = _T_2183 | _T_2184;
  assign _T_2195 = _T_2194 | _T_2185;
  assign _T_2196 = _T_2195 | _T_2186;
  assign _T_2197 = _T_2196 | _T_2187;
  assign _T_2198 = _T_2197 | _T_2188;
  assign _T_2199 = _T_2198 | _T_2189;
  assign _T_2200 = _T_2199 | _T_2190;
  assign _T_2201 = _T_2200 | _T_2191;
  assign _T_2202 = _T_2201 | _T_2192;
  assign _T_2203 = _T_2202 | _T_2193;
  assign _T_2205 = _T_2203 ? io_badaddr : 32'h0;
  assign _T_2213 = causeIsDebugTrigger ? 2'h2 : 2'h1;
  assign _T_2214 = causeIsDebugInt ? 2'h3 : _T_2213;
  assign _T_2215 = reg_singleStepped ? 3'h4 : {{1'd0}, _T_2214};
  assign _GEN_57 = _T_964 ? 1'h1 : reg_debug;
  assign _GEN_58 = _T_964 ? _T_2171 : reg_dpc;
  assign _GEN_59 = _T_964 ? _T_2215 : reg_dcsr_cause;
  assign _GEN_60 = _T_964 ? 2'h3 : reg_dcsr_prv;
  assign _GEN_62 = _T_2071 ? _GEN_57 : reg_debug;
  assign _GEN_63 = _T_2071 ? _GEN_58 : reg_dpc;
  assign _GEN_64 = _T_2071 ? _GEN_59 : reg_dcsr_cause;
  assign _GEN_65 = _T_2071 ? _GEN_60 : reg_dcsr_prv;
  assign _T_2219 = _T_2071 == 1'h0;
  assign _T_2221 = ~ _T_2171;
  assign _T_2222 = reg_misa[2];
  assign _T_2224 = _T_2222 == 1'h0;
  assign _T_2226 = {_T_2224,1'h1};
  assign _GEN_6 = {{30'd0}, _T_2226};
  assign _T_2227 = _T_2221 | _GEN_6;
  assign _T_2228 = ~ _T_2227;
  assign _GEN_71 = {{1'd0}, reg_mstatus_spp};
  assign _GEN_74 = _T_2219 ? _T_2228 : reg_mepc;
  assign _GEN_75 = _T_2219 ? cause : reg_mcause;
  assign _GEN_76 = _T_2219 ? _T_2205 : reg_mbadaddr;
  assign _GEN_77 = _T_2219 ? reg_mstatus_mie : reg_mstatus_mpie;
  assign _GEN_78 = _T_2219 ? 2'h3 : reg_mstatus_mpp;
  assign _GEN_79 = _T_2219 ? 1'h0 : reg_mstatus_mie;
  assign _GEN_81 = exception ? _GEN_62 : reg_debug;
  assign _GEN_82 = exception ? _GEN_63 : reg_dpc;
  assign _GEN_83 = exception ? _GEN_64 : reg_dcsr_cause;
  assign _GEN_84 = exception ? _GEN_65 : reg_dcsr_prv;
  assign _GEN_90 = exception ? _GEN_71 : {{1'd0}, reg_mstatus_spp};
  assign _GEN_92 = exception ? _GEN_74 : reg_mepc;
  assign _GEN_93 = exception ? _GEN_75 : reg_mcause;
  assign _GEN_94 = exception ? _GEN_76 : reg_mbadaddr;
  assign _GEN_95 = exception ? _GEN_77 : reg_mstatus_mpie;
  assign _GEN_96 = exception ? _GEN_78 : reg_mstatus_mpp;
  assign _GEN_97 = exception ? _GEN_79 : reg_mstatus_mie;
  assign _T_2255 = io_rw_addr[10];
  assign _GEN_104 = _T_2255 ? 1'h0 : _GEN_81;
  assign _GEN_105 = _T_2255 ? reg_dpc : tvec;
  assign _T_2264 = _T_2255 == 1'h0;
  assign _GEN_106 = _T_2264 ? reg_mstatus_mpie : _GEN_97;
  assign _GEN_107 = _T_2264 ? 1'h1 : _GEN_95;
  assign _GEN_108 = _T_2264 ? 2'h3 : _GEN_96;
  assign _GEN_110 = _T_2264 ? reg_mepc : _GEN_105;
  assign _GEN_115 = insn_ret ? _GEN_110 : tvec;
  assign _GEN_116 = insn_ret ? _GEN_104 : _GEN_81;
  assign _GEN_117 = insn_ret ? _GEN_106 : _GEN_97;
  assign _GEN_118 = insn_ret ? _GEN_107 : _GEN_95;
  assign _GEN_119 = insn_ret ? _GEN_108 : _GEN_96;
  assign _T_2271 = _T_1249 ? reg_tselect : 1'h0;
  assign _T_2273 = _T_1251 ? _T_1118 : 32'h0;
  assign _T_2275 = _T_1253 ? _GEN_52 : 32'h0;
  assign _T_2283 = _T_1261 ? _T_270 : 64'h0;
  assign _T_2285 = _T_1263 ? _T_257 : 64'h0;
  assign _T_2287 = _T_1265 ? reg_misa : 32'h0;
  assign _T_2289 = _T_1267 ? read_mstatus : 32'h0;
  assign _T_2291 = _T_1269 ? reg_mtvec : 32'h0;
  assign _T_2293 = _T_1271 ? read_mip : 16'h0;
  assign _T_2295 = _T_1273 ? reg_mie : 32'h0;
  assign _T_2297 = _T_1275 ? reg_mscratch : 32'h0;
  assign _T_2299 = _T_1277 ? reg_mepc : 32'h0;
  assign _T_2301 = _T_1279 ? reg_mbadaddr : 32'h0;
  assign _T_2303 = _T_1281 ? reg_mcause : 32'h0;
  assign _T_2305 = _T_1283 ? io_hartid : 1'h0;
  assign _T_2307 = _T_1285 ? _T_1135 : 32'h0;
  assign _T_2309 = _T_1287 ? reg_dpc : 32'h0;
  assign _T_2311 = _T_1289 ? reg_dscratch : 32'h0;
  assign _T_2487 = _T_1465 ? _T_1139 : 32'h0;
  assign _T_2489 = _T_1467 ? _T_1140 : 32'h0;
  assign _T_2491 = _T_1469 ? _T_1178 : 32'h0;
  assign _T_2493 = _T_1471 ? _T_1201 : 32'h0;
  assign _T_2499 = _T_1477 ? reg_pmp_0_addr : 30'h0;
  assign _T_2501 = _T_1479 ? reg_pmp_1_addr : 30'h0;
  assign _T_2503 = _T_1481 ? reg_pmp_2_addr : 30'h0;
  assign _T_2505 = _T_1483 ? reg_pmp_3_addr : 30'h0;
  assign _T_2507 = _T_1485 ? reg_pmp_4_addr : 30'h0;
  assign _T_2509 = _T_1487 ? reg_pmp_5_addr : 30'h0;
  assign _T_2511 = _T_1489 ? reg_pmp_6_addr : 30'h0;
  assign _T_2513 = _T_1491 ? reg_pmp_7_addr : 30'h0;
  assign _GEN_8 = {{31'd0}, _T_2271};
  assign _T_2530 = _GEN_8 | _T_2273;
  assign _T_2531 = _T_2530 | _T_2275;
  assign _GEN_9 = {{32'd0}, _T_2531};
  assign _T_2535 = _GEN_9 | _T_2283;
  assign _T_2536 = _T_2535 | _T_2285;
  assign _GEN_10 = {{32'd0}, _T_2287};
  assign _T_2537 = _T_2536 | _GEN_10;
  assign _GEN_11 = {{32'd0}, _T_2289};
  assign _T_2538 = _T_2537 | _GEN_11;
  assign _GEN_12 = {{32'd0}, _T_2291};
  assign _T_2539 = _T_2538 | _GEN_12;
  assign _GEN_13 = {{48'd0}, _T_2293};
  assign _T_2540 = _T_2539 | _GEN_13;
  assign _GEN_14 = {{32'd0}, _T_2295};
  assign _T_2541 = _T_2540 | _GEN_14;
  assign _GEN_15 = {{32'd0}, _T_2297};
  assign _T_2542 = _T_2541 | _GEN_15;
  assign _GEN_16 = {{32'd0}, _T_2299};
  assign _T_2543 = _T_2542 | _GEN_16;
  assign _GEN_431 = {{32'd0}, _T_2301};
  assign _T_2544 = _T_2543 | _GEN_431;
  assign _GEN_432 = {{32'd0}, _T_2303};
  assign _T_2545 = _T_2544 | _GEN_432;
  assign _GEN_433 = {{63'd0}, _T_2305};
  assign _T_2546 = _T_2545 | _GEN_433;
  assign _GEN_434 = {{32'd0}, _T_2307};
  assign _T_2547 = _T_2546 | _GEN_434;
  assign _GEN_435 = {{32'd0}, _T_2309};
  assign _T_2548 = _T_2547 | _GEN_435;
  assign _GEN_436 = {{32'd0}, _T_2311};
  assign _T_2549 = _T_2548 | _GEN_436;
  assign _GEN_437 = {{32'd0}, _T_2487};
  assign _T_2637 = _T_2549 | _GEN_437;
  assign _GEN_438 = {{32'd0}, _T_2489};
  assign _T_2638 = _T_2637 | _GEN_438;
  assign _GEN_439 = {{32'd0}, _T_2491};
  assign _T_2639 = _T_2638 | _GEN_439;
  assign _GEN_440 = {{32'd0}, _T_2493};
  assign _T_2640 = _T_2639 | _GEN_440;
  assign _GEN_441 = {{34'd0}, _T_2499};
  assign _T_2643 = _T_2640 | _GEN_441;
  assign _GEN_442 = {{34'd0}, _T_2501};
  assign _T_2644 = _T_2643 | _GEN_442;
  assign _GEN_443 = {{34'd0}, _T_2503};
  assign _T_2645 = _T_2644 | _GEN_443;
  assign _GEN_444 = {{34'd0}, _T_2505};
  assign _T_2646 = _T_2645 | _GEN_444;
  assign _GEN_445 = {{34'd0}, _T_2507};
  assign _T_2647 = _T_2646 | _GEN_445;
  assign _GEN_446 = {{34'd0}, _T_2509};
  assign _T_2648 = _T_2647 | _GEN_446;
  assign _GEN_447 = {{34'd0}, _T_2511};
  assign _T_2649 = _T_2648 | _GEN_447;
  assign _GEN_448 = {{34'd0}, _T_2513};
  assign _T_2650 = _T_2649 | _GEN_448;
  assign _T_2667 = io_rw_cmd == 3'h1;
  assign _T_2669 = _T_1512 | _T_2667;
  assign _T_2674 = {{69'd0}, wdata};
  assign _T_2678 = _T_2674[3];
  assign _T_2682 = _T_2674[7];
  assign _GEN_121 = _T_1267 ? _T_2678 : _GEN_117;
  assign _GEN_122 = _T_1267 ? _T_2682 : _GEN_118;
  assign _T_2705 = wdata[5];
  assign _T_2706 = ~ wdata;
  assign _T_2708 = _T_2705 == 1'h0;
  assign _GEN_449 = {{3'd0}, _T_2708};
  assign _T_2709 = _GEN_449 << 3;
  assign _GEN_450 = {{28'd0}, _T_2709};
  assign _T_2710 = _T_2706 | _GEN_450;
  assign _T_2711 = ~ _T_2710;
  assign _T_2712 = _T_2711 & 32'h1005;
  assign _T_2714 = reg_misa & 32'hffffeffa;
  assign _T_2715 = _T_2712 | _T_2714;
  assign _GEN_123 = _T_1265 ? _T_2715 : reg_misa;
  assign _T_2772 = wdata & 32'h888;
  assign _GEN_124 = _T_1273 ? _T_2772 : reg_mie;
  assign _T_2779 = _T_2706 | _GEN_6;
  assign _T_2780 = ~ _T_2779;
  assign _GEN_125 = _T_1277 ? _T_2780 : _GEN_92;
  assign _GEN_126 = _T_1275 ? wdata : reg_mscratch;
  assign _T_2783 = _T_2706 | 32'h2;
  assign _T_2784 = wdata[0];
  assign _T_2787 = _T_2784 ? 6'h3c : 6'h0;
  assign _GEN_453 = {{26'd0}, _T_2787};
  assign _T_2788 = _T_2783 | _GEN_453;
  assign _T_2789 = ~ _T_2788;
  assign _GEN_127 = _T_1269 ? _T_2789 : reg_mtvec;
  assign _T_2791 = wdata & 32'h8000001f;
  assign _GEN_128 = _T_1281 ? _T_2791 : _GEN_93;
  assign _GEN_129 = _T_1279 ? wdata : _GEN_94;
  assign _T_2793 = _T_270[63:32];
  assign _T_2794 = {_T_2793,wdata};
  assign _T_2795 = _T_2794[63:6];
  assign _GEN_130 = _T_1261 ? _T_2794 : {{57'd0}, _T_262};
  assign _GEN_131 = _T_1261 ? _T_2795 : _GEN_36;
  assign _T_2797 = _T_270[31:0];
  assign _T_2798 = {wdata,_T_2797};
  assign _T_2799 = _T_2798[63:6];
  assign _GEN_132 = _T_1465 ? _T_2798 : _GEN_130;
  assign _GEN_133 = _T_1465 ? _T_2799 : _GEN_131;
  assign _T_2800 = _T_257[63:32];
  assign _T_2801 = {_T_2800,wdata};
  assign _T_2802 = _T_2801[63:6];
  assign _GEN_134 = _T_1263 ? _T_2801 : {{57'd0}, _T_249};
  assign _GEN_135 = _T_1263 ? _T_2802 : _GEN_35;
  assign _T_2804 = _T_257[31:0];
  assign _T_2805 = {wdata,_T_2804};
  assign _T_2806 = _T_2805[63:6];
  assign _GEN_136 = _T_1467 ? _T_2805 : _GEN_134;
  assign _GEN_137 = _T_1467 ? _T_2806 : _GEN_135;
  assign _T_2813 = wdata[2];
  assign _T_2819 = wdata[12];
  assign _T_2822 = wdata[15];
  assign _GEN_138 = _T_1285 ? _T_2813 : reg_dcsr_step;
  assign _GEN_139 = _T_1285 ? _T_2822 : reg_dcsr_ebreakm;
  assign _T_2828 = _T_2706 | 32'h1;
  assign _T_2829 = ~ _T_2828;
  assign _GEN_140 = _T_1287 ? _T_2829 : _GEN_82;
  assign _GEN_141 = _T_1289 ? wdata : reg_dscratch;
  assign _T_2832 = _GEN_38 == 1'h0;
  assign _T_2833 = _T_2832 | reg_debug;
  assign _T_2840 = wdata[1];
  assign _T_2846 = wdata[8:7];
  assign _T_2852 = wdata[27];
  assign _T_2854 = _T_2852 & reg_debug;
  assign _GEN_145 = 1'h0 == reg_tselect ? _T_2852 : reg_bp_0_control_dmode;
  assign _GEN_151 = 1'h0 == reg_tselect ? _T_2819 : reg_bp_0_control_action;
  assign _GEN_157 = 1'h0 == reg_tselect ? _T_2846 : reg_bp_0_control_tmatch;
  assign _GEN_167 = 1'h0 == reg_tselect ? _T_2813 : reg_bp_0_control_x;
  assign _GEN_169 = 1'h0 == reg_tselect ? _T_2840 : reg_bp_0_control_w;
  assign _GEN_171 = 1'h0 == reg_tselect ? _T_2784 : reg_bp_0_control_r;
  assign _GEN_173 = 1'h0 == reg_tselect ? _T_2854 : _GEN_145;
  assign _T_2855 = _T_2854 & _T_2819;
  assign _GEN_175 = 1'h0 == reg_tselect ? _T_2855 : _GEN_151;
  assign _GEN_179 = _T_1251 ? _GEN_173 : reg_bp_0_control_dmode;
  assign _GEN_185 = _T_1251 ? _GEN_175 : reg_bp_0_control_action;
  assign _GEN_191 = _T_1251 ? _GEN_157 : reg_bp_0_control_tmatch;
  assign _GEN_201 = _T_1251 ? _GEN_167 : reg_bp_0_control_x;
  assign _GEN_203 = _T_1251 ? _GEN_169 : reg_bp_0_control_w;
  assign _GEN_205 = _T_1251 ? _GEN_171 : reg_bp_0_control_r;
  assign _GEN_207 = 1'h0 == reg_tselect ? wdata : reg_bp_0_address;
  assign _GEN_209 = _T_1253 ? _GEN_207 : reg_bp_0_address;
  assign _GEN_213 = _T_2833 ? _GEN_179 : reg_bp_0_control_dmode;
  assign _GEN_219 = _T_2833 ? _GEN_185 : reg_bp_0_control_action;
  assign _GEN_225 = _T_2833 ? _GEN_191 : reg_bp_0_control_tmatch;
  assign _GEN_235 = _T_2833 ? _GEN_201 : reg_bp_0_control_x;
  assign _GEN_237 = _T_2833 ? _GEN_203 : reg_bp_0_control_w;
  assign _GEN_239 = _T_2833 ? _GEN_205 : reg_bp_0_control_r;
  assign _GEN_241 = _T_2833 ? _GEN_209 : reg_bp_0_address;
  assign _T_2857 = reg_pmp_0_cfg_l == 1'h0;
  assign _T_2858 = _T_1469 & _T_2857;
  assign _T_2864 = wdata[7:0];
  assign _T_2865 = _T_2864[0];
  assign _T_2866 = _T_2864[1];
  assign _T_2867 = _T_2864[2];
  assign _T_2868 = _T_2864[4:3];
  assign _T_2870 = _T_2864[7];
  assign _GEN_243 = _T_2858 ? _T_2870 : reg_pmp_0_cfg_l;
  assign _GEN_245 = _T_2858 ? _T_2868 : reg_pmp_0_cfg_a;
  assign _GEN_246 = _T_2858 ? _T_2867 : reg_pmp_0_cfg_x;
  assign _GEN_247 = _T_2858 ? _T_2866 : reg_pmp_0_cfg_w;
  assign _GEN_248 = _T_2858 ? _T_2865 : reg_pmp_0_cfg_r;
  assign _T_2871 = reg_pmp_1_cfg_a[1];
  assign _T_2872 = reg_pmp_1_cfg_l & _T_2871;
  assign _T_2873 = reg_pmp_0_cfg_l | _T_2872;
  assign _T_2875 = _T_2873 == 1'h0;
  assign _T_2876 = _T_1477 & _T_2875;
  assign _GEN_249 = _T_2876 ? wdata : {{2'd0}, reg_pmp_0_addr};
  assign _T_2878 = reg_pmp_1_cfg_l == 1'h0;
  assign _T_2879 = _T_1469 & _T_2878;
  assign _T_2881 = wdata[31:8];
  assign _T_2885 = _T_2881[7:0];
  assign _T_2886 = _T_2885[0];
  assign _T_2887 = _T_2885[1];
  assign _T_2888 = _T_2885[2];
  assign _T_2889 = _T_2885[4:3];
  assign _T_2891 = _T_2885[7];
  assign _GEN_250 = _T_2879 ? _T_2891 : reg_pmp_1_cfg_l;
  assign _GEN_252 = _T_2879 ? _T_2889 : reg_pmp_1_cfg_a;
  assign _GEN_253 = _T_2879 ? _T_2888 : reg_pmp_1_cfg_x;
  assign _GEN_254 = _T_2879 ? _T_2887 : reg_pmp_1_cfg_w;
  assign _GEN_255 = _T_2879 ? _T_2886 : reg_pmp_1_cfg_r;
  assign _T_2892 = reg_pmp_2_cfg_a[1];
  assign _T_2893 = reg_pmp_2_cfg_l & _T_2892;
  assign _T_2894 = reg_pmp_1_cfg_l | _T_2893;
  assign _T_2896 = _T_2894 == 1'h0;
  assign _T_2897 = _T_1479 & _T_2896;
  assign _GEN_256 = _T_2897 ? wdata : {{2'd0}, reg_pmp_1_addr};
  assign _T_2899 = reg_pmp_2_cfg_l == 1'h0;
  assign _T_2900 = _T_1469 & _T_2899;
  assign _T_2902 = wdata[31:16];
  assign _T_2906 = _T_2902[7:0];
  assign _T_2907 = _T_2906[0];
  assign _T_2908 = _T_2906[1];
  assign _T_2909 = _T_2906[2];
  assign _T_2910 = _T_2906[4:3];
  assign _T_2912 = _T_2906[7];
  assign _GEN_257 = _T_2900 ? _T_2912 : reg_pmp_2_cfg_l;
  assign _GEN_259 = _T_2900 ? _T_2910 : reg_pmp_2_cfg_a;
  assign _GEN_260 = _T_2900 ? _T_2909 : reg_pmp_2_cfg_x;
  assign _GEN_261 = _T_2900 ? _T_2908 : reg_pmp_2_cfg_w;
  assign _GEN_262 = _T_2900 ? _T_2907 : reg_pmp_2_cfg_r;
  assign _T_2913 = reg_pmp_3_cfg_a[1];
  assign _T_2914 = reg_pmp_3_cfg_l & _T_2913;
  assign _T_2915 = reg_pmp_2_cfg_l | _T_2914;
  assign _T_2917 = _T_2915 == 1'h0;
  assign _T_2918 = _T_1481 & _T_2917;
  assign _GEN_263 = _T_2918 ? wdata : {{2'd0}, reg_pmp_2_addr};
  assign _T_2920 = reg_pmp_3_cfg_l == 1'h0;
  assign _T_2921 = _T_1469 & _T_2920;
  assign _T_2923 = wdata[31:24];
  assign _T_2928 = _T_2923[0];
  assign _T_2929 = _T_2923[1];
  assign _T_2930 = _T_2923[2];
  assign _T_2931 = _T_2923[4:3];
  assign _T_2933 = _T_2923[7];
  assign _GEN_264 = _T_2921 ? _T_2933 : reg_pmp_3_cfg_l;
  assign _GEN_266 = _T_2921 ? _T_2931 : reg_pmp_3_cfg_a;
  assign _GEN_267 = _T_2921 ? _T_2930 : reg_pmp_3_cfg_x;
  assign _GEN_268 = _T_2921 ? _T_2929 : reg_pmp_3_cfg_w;
  assign _GEN_269 = _T_2921 ? _T_2928 : reg_pmp_3_cfg_r;
  assign _T_2934 = reg_pmp_4_cfg_a[1];
  assign _T_2935 = reg_pmp_4_cfg_l & _T_2934;
  assign _T_2936 = reg_pmp_3_cfg_l | _T_2935;
  assign _T_2938 = _T_2936 == 1'h0;
  assign _T_2939 = _T_1483 & _T_2938;
  assign _GEN_270 = _T_2939 ? wdata : {{2'd0}, reg_pmp_3_addr};
  assign _T_2941 = reg_pmp_4_cfg_l == 1'h0;
  assign _T_2942 = _T_1471 & _T_2941;
  assign _T_2948 = wdata[7:0];
  assign _T_2949 = _T_2948[0];
  assign _T_2950 = _T_2948[1];
  assign _T_2951 = _T_2948[2];
  assign _T_2952 = _T_2948[4:3];
  assign _T_2954 = _T_2948[7];
  assign _GEN_271 = _T_2942 ? _T_2954 : reg_pmp_4_cfg_l;
  assign _GEN_273 = _T_2942 ? _T_2952 : reg_pmp_4_cfg_a;
  assign _GEN_274 = _T_2942 ? _T_2951 : reg_pmp_4_cfg_x;
  assign _GEN_275 = _T_2942 ? _T_2950 : reg_pmp_4_cfg_w;
  assign _GEN_276 = _T_2942 ? _T_2949 : reg_pmp_4_cfg_r;
  assign _T_2955 = reg_pmp_5_cfg_a[1];
  assign _T_2956 = reg_pmp_5_cfg_l & _T_2955;
  assign _T_2957 = reg_pmp_4_cfg_l | _T_2956;
  assign _T_2959 = _T_2957 == 1'h0;
  assign _T_2960 = _T_1485 & _T_2959;
  assign _GEN_277 = _T_2960 ? wdata : {{2'd0}, reg_pmp_4_addr};
  assign _T_2962 = reg_pmp_5_cfg_l == 1'h0;
  assign _T_2963 = _T_1471 & _T_2962;
  assign _T_2969 = _T_2881[7:0];
  assign _T_2970 = _T_2969[0];
  assign _T_2971 = _T_2969[1];
  assign _T_2972 = _T_2969[2];
  assign _T_2973 = _T_2969[4:3];
  assign _T_2975 = _T_2969[7];
  assign _GEN_278 = _T_2963 ? _T_2975 : reg_pmp_5_cfg_l;
  assign _GEN_280 = _T_2963 ? _T_2973 : reg_pmp_5_cfg_a;
  assign _GEN_281 = _T_2963 ? _T_2972 : reg_pmp_5_cfg_x;
  assign _GEN_282 = _T_2963 ? _T_2971 : reg_pmp_5_cfg_w;
  assign _GEN_283 = _T_2963 ? _T_2970 : reg_pmp_5_cfg_r;
  assign _T_2976 = reg_pmp_6_cfg_a[1];
  assign _T_2977 = reg_pmp_6_cfg_l & _T_2976;
  assign _T_2978 = reg_pmp_5_cfg_l | _T_2977;
  assign _T_2980 = _T_2978 == 1'h0;
  assign _T_2981 = _T_1487 & _T_2980;
  assign _GEN_284 = _T_2981 ? wdata : {{2'd0}, reg_pmp_5_addr};
  assign _T_2983 = reg_pmp_6_cfg_l == 1'h0;
  assign _T_2984 = _T_1471 & _T_2983;
  assign _T_2990 = _T_2902[7:0];
  assign _T_2991 = _T_2990[0];
  assign _T_2992 = _T_2990[1];
  assign _T_2993 = _T_2990[2];
  assign _T_2994 = _T_2990[4:3];
  assign _T_2996 = _T_2990[7];
  assign _GEN_285 = _T_2984 ? _T_2996 : reg_pmp_6_cfg_l;
  assign _GEN_287 = _T_2984 ? _T_2994 : reg_pmp_6_cfg_a;
  assign _GEN_288 = _T_2984 ? _T_2993 : reg_pmp_6_cfg_x;
  assign _GEN_289 = _T_2984 ? _T_2992 : reg_pmp_6_cfg_w;
  assign _GEN_290 = _T_2984 ? _T_2991 : reg_pmp_6_cfg_r;
  assign _T_2997 = reg_pmp_7_cfg_a[1];
  assign _T_2998 = reg_pmp_7_cfg_l & _T_2997;
  assign _T_2999 = reg_pmp_6_cfg_l | _T_2998;
  assign _T_3001 = _T_2999 == 1'h0;
  assign _T_3002 = _T_1489 & _T_3001;
  assign _GEN_291 = _T_3002 ? wdata : {{2'd0}, reg_pmp_6_addr};
  assign _T_3004 = reg_pmp_7_cfg_l == 1'h0;
  assign _T_3005 = _T_1471 & _T_3004;
  assign _GEN_292 = _T_3005 ? _T_2933 : reg_pmp_7_cfg_l;
  assign _GEN_294 = _T_3005 ? _T_2931 : reg_pmp_7_cfg_a;
  assign _GEN_295 = _T_3005 ? _T_2930 : reg_pmp_7_cfg_x;
  assign _GEN_296 = _T_3005 ? _T_2929 : reg_pmp_7_cfg_w;
  assign _GEN_297 = _T_3005 ? _T_2928 : reg_pmp_7_cfg_r;
  assign _T_3020 = reg_pmp_7_cfg_l | _T_2998;
  assign _T_3022 = _T_3020 == 1'h0;
  assign _T_3023 = _T_1491 & _T_3022;
  assign _GEN_298 = _T_3023 ? wdata : {{2'd0}, reg_pmp_7_addr};
  assign _GEN_299 = _T_2669 ? _GEN_121 : _GEN_117;
  assign _GEN_300 = _T_2669 ? _GEN_122 : _GEN_118;
  assign _GEN_301 = _T_2669 ? _GEN_123 : reg_misa;
  assign _GEN_302 = _T_2669 ? _GEN_124 : reg_mie;
  assign _GEN_303 = _T_2669 ? _GEN_125 : _GEN_92;
  assign _GEN_304 = _T_2669 ? _GEN_126 : reg_mscratch;
  assign _GEN_305 = _T_2669 ? _GEN_127 : reg_mtvec;
  assign _GEN_306 = _T_2669 ? _GEN_128 : _GEN_93;
  assign _GEN_307 = _T_2669 ? _GEN_129 : _GEN_94;
  assign _GEN_308 = _T_2669 ? _GEN_132 : {{57'd0}, _T_262};
  assign _GEN_309 = _T_2669 ? _GEN_133 : _GEN_36;
  assign _GEN_310 = _T_2669 ? _GEN_136 : {{57'd0}, _T_249};
  assign _GEN_311 = _T_2669 ? _GEN_137 : _GEN_35;
  assign _GEN_312 = _T_2669 ? _GEN_138 : reg_dcsr_step;
  assign _GEN_313 = _T_2669 ? _GEN_139 : reg_dcsr_ebreakm;
  assign _GEN_314 = _T_2669 ? _GEN_140 : _GEN_82;
  assign _GEN_315 = _T_2669 ? _GEN_141 : reg_dscratch;
  assign _GEN_319 = _T_2669 ? _GEN_213 : reg_bp_0_control_dmode;
  assign _GEN_325 = _T_2669 ? _GEN_219 : reg_bp_0_control_action;
  assign _GEN_331 = _T_2669 ? _GEN_225 : reg_bp_0_control_tmatch;
  assign _GEN_341 = _T_2669 ? _GEN_235 : reg_bp_0_control_x;
  assign _GEN_343 = _T_2669 ? _GEN_237 : reg_bp_0_control_w;
  assign _GEN_345 = _T_2669 ? _GEN_239 : reg_bp_0_control_r;
  assign _GEN_347 = _T_2669 ? _GEN_241 : reg_bp_0_address;
  assign _GEN_349 = _T_2669 ? _GEN_243 : reg_pmp_0_cfg_l;
  assign _GEN_351 = _T_2669 ? _GEN_245 : reg_pmp_0_cfg_a;
  assign _GEN_352 = _T_2669 ? _GEN_246 : reg_pmp_0_cfg_x;
  assign _GEN_353 = _T_2669 ? _GEN_247 : reg_pmp_0_cfg_w;
  assign _GEN_354 = _T_2669 ? _GEN_248 : reg_pmp_0_cfg_r;
  assign _GEN_355 = _T_2669 ? _GEN_249 : {{2'd0}, reg_pmp_0_addr};
  assign _GEN_356 = _T_2669 ? _GEN_250 : reg_pmp_1_cfg_l;
  assign _GEN_358 = _T_2669 ? _GEN_252 : reg_pmp_1_cfg_a;
  assign _GEN_359 = _T_2669 ? _GEN_253 : reg_pmp_1_cfg_x;
  assign _GEN_360 = _T_2669 ? _GEN_254 : reg_pmp_1_cfg_w;
  assign _GEN_361 = _T_2669 ? _GEN_255 : reg_pmp_1_cfg_r;
  assign _GEN_362 = _T_2669 ? _GEN_256 : {{2'd0}, reg_pmp_1_addr};
  assign _GEN_363 = _T_2669 ? _GEN_257 : reg_pmp_2_cfg_l;
  assign _GEN_365 = _T_2669 ? _GEN_259 : reg_pmp_2_cfg_a;
  assign _GEN_366 = _T_2669 ? _GEN_260 : reg_pmp_2_cfg_x;
  assign _GEN_367 = _T_2669 ? _GEN_261 : reg_pmp_2_cfg_w;
  assign _GEN_368 = _T_2669 ? _GEN_262 : reg_pmp_2_cfg_r;
  assign _GEN_369 = _T_2669 ? _GEN_263 : {{2'd0}, reg_pmp_2_addr};
  assign _GEN_370 = _T_2669 ? _GEN_264 : reg_pmp_3_cfg_l;
  assign _GEN_372 = _T_2669 ? _GEN_266 : reg_pmp_3_cfg_a;
  assign _GEN_373 = _T_2669 ? _GEN_267 : reg_pmp_3_cfg_x;
  assign _GEN_374 = _T_2669 ? _GEN_268 : reg_pmp_3_cfg_w;
  assign _GEN_375 = _T_2669 ? _GEN_269 : reg_pmp_3_cfg_r;
  assign _GEN_376 = _T_2669 ? _GEN_270 : {{2'd0}, reg_pmp_3_addr};
  assign _GEN_377 = _T_2669 ? _GEN_271 : reg_pmp_4_cfg_l;
  assign _GEN_379 = _T_2669 ? _GEN_273 : reg_pmp_4_cfg_a;
  assign _GEN_380 = _T_2669 ? _GEN_274 : reg_pmp_4_cfg_x;
  assign _GEN_381 = _T_2669 ? _GEN_275 : reg_pmp_4_cfg_w;
  assign _GEN_382 = _T_2669 ? _GEN_276 : reg_pmp_4_cfg_r;
  assign _GEN_383 = _T_2669 ? _GEN_277 : {{2'd0}, reg_pmp_4_addr};
  assign _GEN_384 = _T_2669 ? _GEN_278 : reg_pmp_5_cfg_l;
  assign _GEN_386 = _T_2669 ? _GEN_280 : reg_pmp_5_cfg_a;
  assign _GEN_387 = _T_2669 ? _GEN_281 : reg_pmp_5_cfg_x;
  assign _GEN_388 = _T_2669 ? _GEN_282 : reg_pmp_5_cfg_w;
  assign _GEN_389 = _T_2669 ? _GEN_283 : reg_pmp_5_cfg_r;
  assign _GEN_390 = _T_2669 ? _GEN_284 : {{2'd0}, reg_pmp_5_addr};
  assign _GEN_391 = _T_2669 ? _GEN_285 : reg_pmp_6_cfg_l;
  assign _GEN_393 = _T_2669 ? _GEN_287 : reg_pmp_6_cfg_a;
  assign _GEN_394 = _T_2669 ? _GEN_288 : reg_pmp_6_cfg_x;
  assign _GEN_395 = _T_2669 ? _GEN_289 : reg_pmp_6_cfg_w;
  assign _GEN_396 = _T_2669 ? _GEN_290 : reg_pmp_6_cfg_r;
  assign _GEN_397 = _T_2669 ? _GEN_291 : {{2'd0}, reg_pmp_6_addr};
  assign _GEN_398 = _T_2669 ? _GEN_292 : reg_pmp_7_cfg_l;
  assign _GEN_400 = _T_2669 ? _GEN_294 : reg_pmp_7_cfg_a;
  assign _GEN_401 = _T_2669 ? _GEN_295 : reg_pmp_7_cfg_x;
  assign _GEN_402 = _T_2669 ? _GEN_296 : reg_pmp_7_cfg_w;
  assign _GEN_403 = _T_2669 ? _GEN_297 : reg_pmp_7_cfg_r;
  assign _GEN_404 = _T_2669 ? _GEN_298 : {{2'd0}, reg_pmp_7_addr};
  assign _GEN_405 = reset ? 1'h0 : _GEN_325;
  assign _GEN_406 = reset ? 1'h0 : _GEN_319;
  assign _GEN_407 = reset ? 1'h0 : _GEN_345;
  assign _GEN_408 = reset ? 1'h0 : _GEN_343;
  assign _GEN_409 = reset ? 1'h0 : _GEN_341;
  assign _GEN_415 = reset ? 2'h0 : _GEN_351;
  assign _GEN_416 = reset ? 1'h0 : _GEN_349;
  assign _GEN_417 = reset ? 2'h0 : _GEN_358;
  assign _GEN_418 = reset ? 1'h0 : _GEN_356;
  assign _GEN_419 = reset ? 2'h0 : _GEN_365;
  assign _GEN_420 = reset ? 1'h0 : _GEN_363;
  assign _GEN_421 = reset ? 2'h0 : _GEN_372;
  assign _GEN_422 = reset ? 1'h0 : _GEN_370;
  assign _GEN_423 = reset ? 2'h0 : _GEN_379;
  assign _GEN_424 = reset ? 1'h0 : _GEN_377;
  assign _GEN_425 = reset ? 2'h0 : _GEN_386;
  assign _GEN_426 = reset ? 1'h0 : _GEN_384;
  assign _GEN_427 = reset ? 2'h0 : _GEN_393;
  assign _GEN_428 = reset ? 1'h0 : _GEN_391;
  assign _GEN_429 = reset ? 2'h0 : _GEN_400;
  assign _GEN_430 = reset ? 1'h0 : _GEN_398;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_mstatus_zero2 = _RAND_1[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_mstatus_zero1 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_mstatus_tsr = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_mstatus_tw = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_mstatus_tvm = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_mstatus_mxr = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  reg_mstatus_sum = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  reg_mstatus_mprv = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  reg_mstatus_xs = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  reg_mstatus_fs = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  reg_mstatus_mpp = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  reg_mstatus_hpp = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  reg_mstatus_spp = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  reg_mstatus_mpie = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  reg_mstatus_hpie = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  reg_mstatus_spie = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  reg_mstatus_upie = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  reg_mstatus_mie = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  reg_mstatus_hie = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  reg_mstatus_sie = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  reg_mstatus_uie = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  reg_dcsr_xdebugver = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  reg_dcsr_zero4 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  reg_dcsr_zero3 = _RAND_24[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  reg_dcsr_ebreakm = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  reg_dcsr_ebreakh = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  reg_dcsr_ebreaks = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  reg_dcsr_ebreaku = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  reg_dcsr_zero2 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  reg_dcsr_stopcycle = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  reg_dcsr_stoptime = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  reg_dcsr_cause = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  reg_dcsr_zero1 = _RAND_33[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  reg_dcsr_step = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  reg_dcsr_prv = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  reg_debugint = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  reg_debug = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  reg_dpc = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  reg_dscratch = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  reg_singleStepped = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  reg_tselect = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  reg_bp_0_control_ttype = _RAND_42[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  reg_bp_0_control_dmode = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  reg_bp_0_control_maskmax = _RAND_44[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  reg_bp_0_control_reserved = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  reg_bp_0_control_action = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  reg_bp_0_control_chain = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  reg_bp_0_control_zero = _RAND_48[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  reg_bp_0_control_tmatch = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  reg_bp_0_control_m = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  reg_bp_0_control_h = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  reg_bp_0_control_s = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  reg_bp_0_control_u = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  reg_bp_0_control_x = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  reg_bp_0_control_w = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  reg_bp_0_control_r = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  reg_bp_0_address = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  reg_bp_1_control_ttype = _RAND_58[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  reg_bp_1_control_dmode = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  reg_bp_1_control_maskmax = _RAND_60[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  reg_bp_1_control_reserved = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  reg_bp_1_control_action = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  reg_bp_1_control_chain = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  reg_bp_1_control_zero = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  reg_bp_1_control_tmatch = _RAND_65[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  reg_bp_1_control_m = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  reg_bp_1_control_h = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  reg_bp_1_control_s = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  reg_bp_1_control_u = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  reg_bp_1_control_x = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  reg_bp_1_control_w = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  reg_bp_1_control_r = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  reg_bp_1_address = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  reg_pmp_0_cfg_l = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  reg_pmp_0_cfg_res = _RAND_75[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  reg_pmp_0_cfg_a = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  reg_pmp_0_cfg_x = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  reg_pmp_0_cfg_w = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  reg_pmp_0_cfg_r = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  reg_pmp_0_addr = _RAND_80[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  reg_pmp_1_cfg_l = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  reg_pmp_1_cfg_res = _RAND_82[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  reg_pmp_1_cfg_a = _RAND_83[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  reg_pmp_1_cfg_x = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  reg_pmp_1_cfg_w = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  reg_pmp_1_cfg_r = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  reg_pmp_1_addr = _RAND_87[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  reg_pmp_2_cfg_l = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  reg_pmp_2_cfg_res = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  reg_pmp_2_cfg_a = _RAND_90[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  reg_pmp_2_cfg_x = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  reg_pmp_2_cfg_w = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  reg_pmp_2_cfg_r = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  reg_pmp_2_addr = _RAND_94[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  reg_pmp_3_cfg_l = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  reg_pmp_3_cfg_res = _RAND_96[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  reg_pmp_3_cfg_a = _RAND_97[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  reg_pmp_3_cfg_x = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  reg_pmp_3_cfg_w = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  reg_pmp_3_cfg_r = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  reg_pmp_3_addr = _RAND_101[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  reg_pmp_4_cfg_l = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  reg_pmp_4_cfg_res = _RAND_103[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  reg_pmp_4_cfg_a = _RAND_104[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  reg_pmp_4_cfg_x = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  reg_pmp_4_cfg_w = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  reg_pmp_4_cfg_r = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  reg_pmp_4_addr = _RAND_108[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  reg_pmp_5_cfg_l = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  reg_pmp_5_cfg_res = _RAND_110[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  reg_pmp_5_cfg_a = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  reg_pmp_5_cfg_x = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  reg_pmp_5_cfg_w = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  reg_pmp_5_cfg_r = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  reg_pmp_5_addr = _RAND_115[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  reg_pmp_6_cfg_l = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  reg_pmp_6_cfg_res = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  reg_pmp_6_cfg_a = _RAND_118[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  reg_pmp_6_cfg_x = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  reg_pmp_6_cfg_w = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  reg_pmp_6_cfg_r = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  reg_pmp_6_addr = _RAND_122[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  reg_pmp_7_cfg_l = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  reg_pmp_7_cfg_res = _RAND_124[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  reg_pmp_7_cfg_a = _RAND_125[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  reg_pmp_7_cfg_x = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  reg_pmp_7_cfg_w = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  reg_pmp_7_cfg_r = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  reg_pmp_7_addr = _RAND_129[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  reg_mie = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  reg_mideleg = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  reg_mip_zero2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  reg_mip_debug = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  reg_mip_zero1 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  reg_mip_meip = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  reg_mip_heip = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  reg_mip_seip = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  reg_mip_ueip = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  reg_mip_mtip = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  reg_mip_htip = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  reg_mip_stip = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  reg_mip_utip = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  reg_mip_msip = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  reg_mip_hsip = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  reg_mip_ssip = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  reg_mip_usip = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  reg_mepc = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  reg_mcause = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  reg_mbadaddr = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  reg_mscratch = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  reg_mtvec = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  reg_mcounteren = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  reg_sptbr_ppn = _RAND_153[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  reg_wfi = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_248 = _RAND_155[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {2{$random}};
  _T_252 = _RAND_156[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_261 = _RAND_157[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {2{$random}};
  _T_265 = _RAND_158[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  reg_misa = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_2116 = _RAND_160[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      reg_mstatus_prv <= 2'h3;
    end
    if (reset) begin
      reg_mstatus_zero2 <= 27'h0;
    end
    if (reset) begin
      reg_mstatus_zero1 <= 8'h0;
    end
    if (reset) begin
      reg_mstatus_tsr <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_tw <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_tvm <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_mxr <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_sum <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_mprv <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_xs <= 2'h0;
    end
    if (reset) begin
      reg_mstatus_fs <= 2'h0;
    end
    if (reset) begin
      reg_mstatus_mpp <= 2'h3;
    end else begin
      if (insn_ret) begin
        if (_T_2264) begin
          reg_mstatus_mpp <= 2'h3;
        end else begin
          if (exception) begin
            if (_T_2219) begin
              reg_mstatus_mpp <= 2'h3;
            end
          end
        end
      end else begin
        if (exception) begin
          if (_T_2219) begin
            reg_mstatus_mpp <= 2'h3;
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_hpp <= 2'h0;
    end
    if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_90[0];
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1267) begin
          reg_mstatus_mpie <= _T_2682;
        end else begin
          if (insn_ret) begin
            if (_T_2264) begin
              reg_mstatus_mpie <= 1'h1;
            end else begin
              if (exception) begin
                if (_T_2219) begin
                  reg_mstatus_mpie <= reg_mstatus_mie;
                end
              end
            end
          end else begin
            if (exception) begin
              if (_T_2219) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2264) begin
            reg_mstatus_mpie <= 1'h1;
          end else begin
            if (exception) begin
              if (_T_2219) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end else begin
          if (exception) begin
            if (_T_2219) begin
              reg_mstatus_mpie <= reg_mstatus_mie;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_hpie <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_spie <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_upie <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1267) begin
          reg_mstatus_mie <= _T_2678;
        end else begin
          if (insn_ret) begin
            if (_T_2264) begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end else begin
              if (exception) begin
                if (_T_2219) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            if (exception) begin
              if (_T_2219) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_2264) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end else begin
            if (exception) begin
              if (_T_2219) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end else begin
          if (exception) begin
            if (_T_2219) begin
              reg_mstatus_mie <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_hie <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_sie <= 1'h0;
    end
    if (reset) begin
      reg_mstatus_uie <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_xdebugver <= 2'h1;
    end
    if (reset) begin
      reg_dcsr_zero4 <= 2'h0;
    end
    if (reset) begin
      reg_dcsr_zero3 <= 12'h0;
    end
    if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1285) begin
          reg_dcsr_ebreakm <= _T_2822;
        end
      end
    end
    if (reset) begin
      reg_dcsr_ebreakh <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_ebreaks <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_ebreaku <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_zero2 <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_stopcycle <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_stoptime <= 1'h0;
    end
    if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else begin
      if (exception) begin
        if (_T_2071) begin
          if (_T_964) begin
            if (reg_singleStepped) begin
              reg_dcsr_cause <= 3'h4;
            end else begin
              reg_dcsr_cause <= {{1'd0}, _T_2214};
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_zero1 <= 3'h0;
    end
    if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1285) begin
          reg_dcsr_step <= _T_2813;
        end
      end
    end
    if (reset) begin
      reg_dcsr_prv <= 2'h3;
    end else begin
      if (exception) begin
        if (_T_2071) begin
          if (_T_964) begin
            reg_dcsr_prv <= 2'h3;
          end
        end
      end
    end
    reg_debugint <= io_interrupts_debug;
    if (reset) begin
      reg_debug <= 1'h0;
    end else begin
      if (insn_ret) begin
        if (_T_2255) begin
          reg_debug <= 1'h0;
        end else begin
          if (exception) begin
            if (_T_2071) begin
              if (_T_964) begin
                reg_debug <= 1'h1;
              end
            end
          end
        end
      end else begin
        if (exception) begin
          if (_T_2071) begin
            if (_T_964) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end
    end
    if (_T_2669) begin
      if (_T_1287) begin
        reg_dpc <= _T_2829;
      end else begin
        if (exception) begin
          if (_T_2071) begin
            if (_T_964) begin
              reg_dpc <= _T_2171;
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (_T_2071) begin
          if (_T_964) begin
            reg_dpc <= _T_2171;
          end
        end
      end
    end
    if (_T_2669) begin
      if (_T_1289) begin
        reg_dscratch <= wdata;
      end
    end
    if (_T_967) begin
      reg_singleStepped <= 1'h0;
    end else begin
      if (_T_2147) begin
        reg_singleStepped <= 1'h1;
      end
    end
    reg_tselect <= 1'h0;
    reg_bp_0_control_ttype <= 4'h2;
    if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2833) begin
          if (_T_1251) begin
            if (1'h0 == reg_tselect) begin
              reg_bp_0_control_dmode <= _T_2854;
            end else begin
              if (1'h0 == reg_tselect) begin
                reg_bp_0_control_dmode <= _T_2852;
              end
            end
          end
        end
      end
    end
    reg_bp_0_control_maskmax <= 6'h4;
    reg_bp_0_control_reserved <= 8'h0;
    if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2833) begin
          if (_T_1251) begin
            if (1'h0 == reg_tselect) begin
              reg_bp_0_control_action <= _T_2855;
            end else begin
              if (1'h0 == reg_tselect) begin
                reg_bp_0_control_action <= _T_2819;
              end
            end
          end
        end
      end
    end
    reg_bp_0_control_chain <= 1'h0;
    reg_bp_0_control_zero <= 2'h0;
    if (_T_2669) begin
      if (_T_2833) begin
        if (_T_1251) begin
          if (1'h0 == reg_tselect) begin
            reg_bp_0_control_tmatch <= _T_2846;
          end
        end
      end
    end
    reg_bp_0_control_m <= 1'h1;
    reg_bp_0_control_h <= 1'h0;
    reg_bp_0_control_s <= 1'h0;
    reg_bp_0_control_u <= 1'h0;
    if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2833) begin
          if (_T_1251) begin
            if (1'h0 == reg_tselect) begin
              reg_bp_0_control_x <= _T_2813;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2833) begin
          if (_T_1251) begin
            if (1'h0 == reg_tselect) begin
              reg_bp_0_control_w <= _T_2840;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2833) begin
          if (_T_1251) begin
            if (1'h0 == reg_tselect) begin
              reg_bp_0_control_r <= _T_2784;
            end
          end
        end
      end
    end
    if (_T_2669) begin
      if (_T_2833) begin
        if (_T_1253) begin
          if (1'h0 == reg_tselect) begin
            reg_bp_0_address <= wdata;
          end
        end
      end
    end
    reg_bp_1_control_ttype <= 4'h0;
    reg_bp_1_control_dmode <= 1'h0;
    reg_bp_1_control_maskmax <= 6'h0;
    reg_bp_1_control_reserved <= 8'h0;
    reg_bp_1_control_action <= 1'h0;
    reg_bp_1_control_chain <= 1'h0;
    reg_bp_1_control_zero <= 2'h0;
    reg_bp_1_control_tmatch <= 2'h0;
    reg_bp_1_control_m <= 1'h0;
    reg_bp_1_control_h <= 1'h0;
    reg_bp_1_control_s <= 1'h0;
    reg_bp_1_control_u <= 1'h0;
    reg_bp_1_control_x <= 1'h0;
    reg_bp_1_control_w <= 1'h0;
    reg_bp_1_control_r <= 1'h0;
    reg_bp_1_address <= 32'h0;
    if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2858) begin
          reg_pmp_0_cfg_l <= _T_2870;
        end
      end
    end
    reg_pmp_0_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2858) begin
          reg_pmp_0_cfg_a <= _T_2868;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2858) begin
        reg_pmp_0_cfg_x <= _T_2867;
      end
    end
    if (_T_2669) begin
      if (_T_2858) begin
        reg_pmp_0_cfg_w <= _T_2866;
      end
    end
    if (_T_2669) begin
      if (_T_2858) begin
        reg_pmp_0_cfg_r <= _T_2865;
      end
    end
    reg_pmp_0_addr <= _GEN_355[29:0];
    if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2879) begin
          reg_pmp_1_cfg_l <= _T_2891;
        end
      end
    end
    reg_pmp_1_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2879) begin
          reg_pmp_1_cfg_a <= _T_2889;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2879) begin
        reg_pmp_1_cfg_x <= _T_2888;
      end
    end
    if (_T_2669) begin
      if (_T_2879) begin
        reg_pmp_1_cfg_w <= _T_2887;
      end
    end
    if (_T_2669) begin
      if (_T_2879) begin
        reg_pmp_1_cfg_r <= _T_2886;
      end
    end
    reg_pmp_1_addr <= _GEN_362[29:0];
    if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2900) begin
          reg_pmp_2_cfg_l <= _T_2912;
        end
      end
    end
    reg_pmp_2_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2900) begin
          reg_pmp_2_cfg_a <= _T_2910;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2900) begin
        reg_pmp_2_cfg_x <= _T_2909;
      end
    end
    if (_T_2669) begin
      if (_T_2900) begin
        reg_pmp_2_cfg_w <= _T_2908;
      end
    end
    if (_T_2669) begin
      if (_T_2900) begin
        reg_pmp_2_cfg_r <= _T_2907;
      end
    end
    reg_pmp_2_addr <= _GEN_369[29:0];
    if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2921) begin
          reg_pmp_3_cfg_l <= _T_2933;
        end
      end
    end
    reg_pmp_3_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2921) begin
          reg_pmp_3_cfg_a <= _T_2931;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2921) begin
        reg_pmp_3_cfg_x <= _T_2930;
      end
    end
    if (_T_2669) begin
      if (_T_2921) begin
        reg_pmp_3_cfg_w <= _T_2929;
      end
    end
    if (_T_2669) begin
      if (_T_2921) begin
        reg_pmp_3_cfg_r <= _T_2928;
      end
    end
    reg_pmp_3_addr <= _GEN_376[29:0];
    if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2942) begin
          reg_pmp_4_cfg_l <= _T_2954;
        end
      end
    end
    reg_pmp_4_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2942) begin
          reg_pmp_4_cfg_a <= _T_2952;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2942) begin
        reg_pmp_4_cfg_x <= _T_2951;
      end
    end
    if (_T_2669) begin
      if (_T_2942) begin
        reg_pmp_4_cfg_w <= _T_2950;
      end
    end
    if (_T_2669) begin
      if (_T_2942) begin
        reg_pmp_4_cfg_r <= _T_2949;
      end
    end
    reg_pmp_4_addr <= _GEN_383[29:0];
    if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2963) begin
          reg_pmp_5_cfg_l <= _T_2975;
        end
      end
    end
    reg_pmp_5_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2963) begin
          reg_pmp_5_cfg_a <= _T_2973;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2963) begin
        reg_pmp_5_cfg_x <= _T_2972;
      end
    end
    if (_T_2669) begin
      if (_T_2963) begin
        reg_pmp_5_cfg_w <= _T_2971;
      end
    end
    if (_T_2669) begin
      if (_T_2963) begin
        reg_pmp_5_cfg_r <= _T_2970;
      end
    end
    reg_pmp_5_addr <= _GEN_390[29:0];
    if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2984) begin
          reg_pmp_6_cfg_l <= _T_2996;
        end
      end
    end
    reg_pmp_6_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_2984) begin
          reg_pmp_6_cfg_a <= _T_2994;
        end
      end
    end
    if (_T_2669) begin
      if (_T_2984) begin
        reg_pmp_6_cfg_x <= _T_2993;
      end
    end
    if (_T_2669) begin
      if (_T_2984) begin
        reg_pmp_6_cfg_w <= _T_2992;
      end
    end
    if (_T_2669) begin
      if (_T_2984) begin
        reg_pmp_6_cfg_r <= _T_2991;
      end
    end
    reg_pmp_6_addr <= _GEN_397[29:0];
    if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else begin
      if (_T_2669) begin
        if (_T_3005) begin
          reg_pmp_7_cfg_l <= _T_2933;
        end
      end
    end
    reg_pmp_7_cfg_res <= 2'h0;
    if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else begin
      if (_T_2669) begin
        if (_T_3005) begin
          reg_pmp_7_cfg_a <= _T_2931;
        end
      end
    end
    if (_T_2669) begin
      if (_T_3005) begin
        reg_pmp_7_cfg_x <= _T_2930;
      end
    end
    if (_T_2669) begin
      if (_T_3005) begin
        reg_pmp_7_cfg_w <= _T_2929;
      end
    end
    if (_T_2669) begin
      if (_T_3005) begin
        reg_pmp_7_cfg_r <= _T_2928;
      end
    end
    reg_pmp_7_addr <= _GEN_404[29:0];
    if (_T_2669) begin
      if (_T_1273) begin
        reg_mie <= _T_2772;
      end
    end
    reg_mideleg <= 32'h0;
    reg_mip_meip <= io_interrupts_meip;
    reg_mip_mtip <= io_interrupts_mtip;
    reg_mip_msip <= io_interrupts_msip;
    if (_T_2669) begin
      if (_T_1277) begin
        reg_mepc <= _T_2780;
      end else begin
        if (exception) begin
          if (_T_2219) begin
            reg_mepc <= _T_2228;
          end
        end
      end
    end else begin
      if (exception) begin
        if (_T_2219) begin
          reg_mepc <= _T_2228;
        end
      end
    end
    if (_T_2669) begin
      if (_T_1281) begin
        reg_mcause <= _T_2791;
      end else begin
        if (exception) begin
          if (_T_2219) begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_2047};
            end else begin
              if (insn_break) begin
                reg_mcause <= 32'h3;
              end else begin
                reg_mcause <= io_cause;
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (_T_2219) begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_2047};
          end else begin
            if (insn_break) begin
              reg_mcause <= 32'h3;
            end else begin
              reg_mcause <= io_cause;
            end
          end
        end
      end
    end
    if (_T_2669) begin
      if (_T_1279) begin
        reg_mbadaddr <= wdata;
      end else begin
        if (exception) begin
          if (_T_2219) begin
            if (_T_2203) begin
              reg_mbadaddr <= io_badaddr;
            end else begin
              reg_mbadaddr <= 32'h0;
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (_T_2219) begin
          if (_T_2203) begin
            reg_mbadaddr <= io_badaddr;
          end else begin
            reg_mbadaddr <= 32'h0;
          end
        end
      end
    end
    if (_T_2669) begin
      if (_T_1275) begin
        reg_mscratch <= wdata;
      end
    end
    if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1269) begin
          reg_mtvec <= _T_2789;
        end
      end
    end
    reg_mcounteren <= 32'h0;
    if (reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if (_T_2136) begin
        reg_wfi <= 1'h0;
      end else begin
        if (_T_2131) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_248 <= 6'h0;
    end else begin
      _T_248 <= _GEN_310[5:0];
    end
    if (reset) begin
      _T_252 <= 58'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1467) begin
          _T_252 <= _T_2806;
        end else begin
          if (_T_1263) begin
            _T_252 <= _T_2802;
          end else begin
            if (_T_253) begin
              _T_252 <= _T_256;
            end
          end
        end
      end else begin
        if (_T_253) begin
          _T_252 <= _T_256;
        end
      end
    end
    if (reset) begin
      _T_261 <= 6'h0;
    end else begin
      _T_261 <= _GEN_308[5:0];
    end
    if (reset) begin
      _T_265 <= 58'h0;
    end else begin
      if (_T_2669) begin
        if (_T_1465) begin
          _T_265 <= _T_2799;
        end else begin
          if (_T_1261) begin
            _T_265 <= _T_2795;
          end else begin
            if (_T_266) begin
              _T_265 <= _T_269;
            end
          end
        end
      end else begin
        if (_T_266) begin
          _T_265 <= _T_269;
        end
      end
    end
    if (reset) begin
      reg_misa <= 32'h40001105;
    end else begin
      if (_T_2669) begin
        if (_T_1265) begin
          reg_misa <= _T_2715;
        end
      end
    end
    if (_T_2113) begin
      _T_2116 <= reg_mstatus_mpp;
    end else begin
      _T_2116 <= reg_mstatus_prv;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2125) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:498 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2145) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:502 assert(!reg_wfi || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2145) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:506 assert(!io.singleStep || io.retire <= UInt(1))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2167) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:507 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2167) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BreakpointUnit(
  input         io_status_debug,
  input  [1:0]  io_status_prv,
  input         io_bp_0_control_action,
  input         io_bp_0_control_chain,
  input  [1:0]  io_bp_0_control_tmatch,
  input         io_bp_0_control_m,
  input         io_bp_0_control_h,
  input         io_bp_0_control_s,
  input         io_bp_0_control_u,
  input         io_bp_0_control_x,
  input         io_bp_0_control_w,
  input         io_bp_0_control_r,
  input  [31:0] io_bp_0_address,
  input  [31:0] io_pc,
  input  [31:0] io_ea,
  output        io_xcpt_if,
  output        io_xcpt_ld,
  output        io_xcpt_st,
  output        io_debug_if,
  output        io_debug_ld,
  output        io_debug_st
);
  wire  _T_27;
  wire [1:0] _T_28;
  wire [1:0] _T_29;
  wire [3:0] _T_30;
  wire [3:0] _T_31;
  wire  _T_32;
  wire  _T_33;
  wire  _T_35;
  wire  _T_36;
  wire  _T_37;
  wire  _T_38;
  wire  _T_39;
  wire [31:0] _T_40;
  wire  _T_42;
  wire  _T_43;
  wire  _T_44;
  wire  _T_45;
  wire  _T_46;
  wire  _T_47;
  wire [1:0] _T_48;
  wire [1:0] _T_49;
  wire [3:0] _T_50;
  wire [31:0] _GEN_6;
  wire [31:0] _T_51;
  wire [31:0] _T_52;
  wire [31:0] _T_63;
  wire  _T_64;
  wire  _T_65;
  wire  _T_66;
  wire  _T_68;
  wire  _T_99;
  wire  _T_101;
  wire  _T_103;
  wire  _T_105;
  wire [31:0] _T_106;
  wire [31:0] _T_117;
  wire  _T_130;
  wire  _T_131;
  wire  _T_132;
  wire  _T_134;
  wire  _T_135;
  wire  _T_137;
  wire  _GEN_0;
  wire  _GEN_1;
  wire  _T_138;
  wire  _GEN_2;
  wire  _GEN_3;
  wire  _T_141;
  wire  _GEN_4;
  wire  _GEN_5;
  assign io_xcpt_if = _GEN_4;
  assign io_xcpt_ld = _GEN_0;
  assign io_xcpt_st = _GEN_2;
  assign io_debug_if = _GEN_5;
  assign io_debug_ld = _GEN_1;
  assign io_debug_st = _GEN_3;
  assign _T_27 = io_status_debug == 1'h0;
  assign _T_28 = {io_bp_0_control_s,io_bp_0_control_u};
  assign _T_29 = {io_bp_0_control_m,io_bp_0_control_h};
  assign _T_30 = {_T_29,_T_28};
  assign _T_31 = _T_30 >> io_status_prv;
  assign _T_32 = _T_31[0];
  assign _T_33 = _T_27 & _T_32;
  assign _T_35 = _T_33 & io_bp_0_control_r;
  assign _T_36 = io_bp_0_control_tmatch[1];
  assign _T_37 = io_ea >= io_bp_0_address;
  assign _T_38 = io_bp_0_control_tmatch[0];
  assign _T_39 = _T_37 ^ _T_38;
  assign _T_40 = ~ io_ea;
  assign _T_42 = io_bp_0_address[0];
  assign _T_43 = _T_38 & _T_42;
  assign _T_44 = io_bp_0_address[1];
  assign _T_45 = _T_43 & _T_44;
  assign _T_46 = io_bp_0_address[2];
  assign _T_47 = _T_45 & _T_46;
  assign _T_48 = {_T_43,_T_38};
  assign _T_49 = {_T_47,_T_45};
  assign _T_50 = {_T_49,_T_48};
  assign _GEN_6 = {{28'd0}, _T_50};
  assign _T_51 = _T_40 | _GEN_6;
  assign _T_52 = ~ io_bp_0_address;
  assign _T_63 = _T_52 | _GEN_6;
  assign _T_64 = _T_51 == _T_63;
  assign _T_65 = _T_36 ? _T_39 : _T_64;
  assign _T_66 = _T_35 & _T_65;
  assign _T_68 = _T_33 & io_bp_0_control_w;
  assign _T_99 = _T_68 & _T_65;
  assign _T_101 = _T_33 & io_bp_0_control_x;
  assign _T_103 = io_pc >= io_bp_0_address;
  assign _T_105 = _T_103 ^ _T_38;
  assign _T_106 = ~ io_pc;
  assign _T_117 = _T_106 | _GEN_6;
  assign _T_130 = _T_117 == _T_63;
  assign _T_131 = _T_36 ? _T_105 : _T_130;
  assign _T_132 = _T_101 & _T_131;
  assign _T_134 = io_bp_0_control_chain == 1'h0;
  assign _T_135 = _T_134 & _T_66;
  assign _T_137 = io_bp_0_control_action == 1'h0;
  assign _GEN_0 = _T_135 ? _T_137 : 1'h0;
  assign _GEN_1 = _T_135 ? io_bp_0_control_action : 1'h0;
  assign _T_138 = _T_134 & _T_99;
  assign _GEN_2 = _T_138 ? _T_137 : 1'h0;
  assign _GEN_3 = _T_138 ? io_bp_0_control_action : 1'h0;
  assign _T_141 = _T_134 & _T_132;
  assign _GEN_4 = _T_141 ? _T_137 : 1'h0;
  assign _GEN_5 = _T_141 ? io_bp_0_control_action : 1'h0;
endmodule
module ALU(
  input  [3:0]  io_fn,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  output [31:0] io_out,
  output [31:0] io_adder_out,
  output        io_cmp_out
);
  wire  _T_9;
  wire [31:0] _T_10;
  wire [31:0] in2_inv;
  wire [31:0] in1_xor_in2;
  wire [32:0] _T_11;
  wire [31:0] _T_12;
  wire [31:0] _GEN_0;
  wire [32:0] _T_14;
  wire [31:0] _T_15;
  wire  _T_16;
  wire  _T_19;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_26;
  wire  _T_29;
  wire  _T_30;
  wire  _T_31;
  wire  _T_32;
  wire [4:0] shamt;
  wire  _T_34;
  wire  _T_36;
  wire  _T_37;
  wire [15:0] _T_42;
  wire [31:0] _T_43;
  wire [15:0] _T_44;
  wire [31:0] _GEN_1;
  wire [31:0] _T_45;
  wire [31:0] _T_47;
  wire [31:0] _T_48;
  wire [23:0] _T_52;
  wire [31:0] _GEN_2;
  wire [31:0] _T_53;
  wire [23:0] _T_54;
  wire [31:0] _GEN_3;
  wire [31:0] _T_55;
  wire [31:0] _T_57;
  wire [31:0] _T_58;
  wire [27:0] _T_62;
  wire [31:0] _GEN_4;
  wire [31:0] _T_63;
  wire [27:0] _T_64;
  wire [31:0] _GEN_5;
  wire [31:0] _T_65;
  wire [31:0] _T_67;
  wire [31:0] _T_68;
  wire [29:0] _T_72;
  wire [31:0] _GEN_6;
  wire [31:0] _T_73;
  wire [29:0] _T_74;
  wire [31:0] _GEN_7;
  wire [31:0] _T_75;
  wire [31:0] _T_77;
  wire [31:0] _T_78;
  wire [30:0] _T_82;
  wire [31:0] _GEN_8;
  wire [31:0] _T_83;
  wire [30:0] _T_84;
  wire [31:0] _GEN_9;
  wire [31:0] _T_85;
  wire [31:0] _T_87;
  wire [31:0] _T_88;
  wire [31:0] shin;
  wire  _T_90;
  wire  _T_91;
  wire [32:0] _T_92;
  wire [32:0] _T_93;
  wire [32:0] _T_94;
  wire [31:0] shout_r;
  wire [15:0] _T_99;
  wire [31:0] _T_100;
  wire [15:0] _T_101;
  wire [31:0] _GEN_10;
  wire [31:0] _T_102;
  wire [31:0] _T_104;
  wire [31:0] _T_105;
  wire [23:0] _T_109;
  wire [31:0] _GEN_11;
  wire [31:0] _T_110;
  wire [23:0] _T_111;
  wire [31:0] _GEN_12;
  wire [31:0] _T_112;
  wire [31:0] _T_114;
  wire [31:0] _T_115;
  wire [27:0] _T_119;
  wire [31:0] _GEN_13;
  wire [31:0] _T_120;
  wire [27:0] _T_121;
  wire [31:0] _GEN_14;
  wire [31:0] _T_122;
  wire [31:0] _T_124;
  wire [31:0] _T_125;
  wire [29:0] _T_129;
  wire [31:0] _GEN_15;
  wire [31:0] _T_130;
  wire [29:0] _T_131;
  wire [31:0] _GEN_16;
  wire [31:0] _T_132;
  wire [31:0] _T_134;
  wire [31:0] _T_135;
  wire [30:0] _T_139;
  wire [31:0] _GEN_17;
  wire [31:0] _T_140;
  wire [30:0] _T_141;
  wire [31:0] _GEN_18;
  wire [31:0] _T_142;
  wire [31:0] _T_144;
  wire [31:0] shout_l;
  wire [31:0] _T_151;
  wire  _T_153;
  wire [31:0] _T_155;
  wire [31:0] shout;
  wire  _T_157;
  wire  _T_159;
  wire  _T_160;
  wire [31:0] _T_162;
  wire  _T_166;
  wire  _T_167;
  wire [31:0] _T_168;
  wire [31:0] _T_170;
  wire [31:0] logic$;
  wire  _T_172;
  wire  _T_174;
  wire  _T_175;
  wire  _T_177;
  wire  _T_178;
  wire  _T_179;
  wire [31:0] _GEN_19;
  wire [31:0] _T_180;
  wire [31:0] shift_logic;
  wire  _T_182;
  wire  _T_184;
  wire  _T_185;
  wire [31:0] out;
  assign io_out = out;
  assign io_adder_out = _T_15;
  assign io_cmp_out = _T_32;
  assign _T_9 = io_fn[3];
  assign _T_10 = ~ io_in2;
  assign in2_inv = _T_9 ? _T_10 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign _T_11 = io_in1 + in2_inv;
  assign _T_12 = _T_11[31:0];
  assign _GEN_0 = {{31'd0}, _T_9};
  assign _T_14 = _T_12 + _GEN_0;
  assign _T_15 = _T_14[31:0];
  assign _T_16 = io_fn[0];
  assign _T_19 = _T_9 == 1'h0;
  assign _T_21 = in1_xor_in2 == 32'h0;
  assign _T_22 = io_in1[31];
  assign _T_23 = io_in2[31];
  assign _T_24 = _T_22 == _T_23;
  assign _T_25 = io_adder_out[31];
  assign _T_26 = io_fn[1];
  assign _T_29 = _T_26 ? _T_23 : _T_22;
  assign _T_30 = _T_24 ? _T_25 : _T_29;
  assign _T_31 = _T_19 ? _T_21 : _T_30;
  assign _T_32 = _T_16 ^ _T_31;
  assign shamt = io_in2[4:0];
  assign _T_34 = io_fn == 4'h5;
  assign _T_36 = io_fn == 4'hb;
  assign _T_37 = _T_34 | _T_36;
  assign _T_42 = io_in1[31:16];
  assign _T_43 = {{16'd0}, _T_42};
  assign _T_44 = io_in1[15:0];
  assign _GEN_1 = {{16'd0}, _T_44};
  assign _T_45 = _GEN_1 << 16;
  assign _T_47 = _T_45 & 32'hffff0000;
  assign _T_48 = _T_43 | _T_47;
  assign _T_52 = _T_48[31:8];
  assign _GEN_2 = {{8'd0}, _T_52};
  assign _T_53 = _GEN_2 & 32'hff00ff;
  assign _T_54 = _T_48[23:0];
  assign _GEN_3 = {{8'd0}, _T_54};
  assign _T_55 = _GEN_3 << 8;
  assign _T_57 = _T_55 & 32'hff00ff00;
  assign _T_58 = _T_53 | _T_57;
  assign _T_62 = _T_58[31:4];
  assign _GEN_4 = {{4'd0}, _T_62};
  assign _T_63 = _GEN_4 & 32'hf0f0f0f;
  assign _T_64 = _T_58[27:0];
  assign _GEN_5 = {{4'd0}, _T_64};
  assign _T_65 = _GEN_5 << 4;
  assign _T_67 = _T_65 & 32'hf0f0f0f0;
  assign _T_68 = _T_63 | _T_67;
  assign _T_72 = _T_68[31:2];
  assign _GEN_6 = {{2'd0}, _T_72};
  assign _T_73 = _GEN_6 & 32'h33333333;
  assign _T_74 = _T_68[29:0];
  assign _GEN_7 = {{2'd0}, _T_74};
  assign _T_75 = _GEN_7 << 2;
  assign _T_77 = _T_75 & 32'hcccccccc;
  assign _T_78 = _T_73 | _T_77;
  assign _T_82 = _T_78[31:1];
  assign _GEN_8 = {{1'd0}, _T_82};
  assign _T_83 = _GEN_8 & 32'h55555555;
  assign _T_84 = _T_78[30:0];
  assign _GEN_9 = {{1'd0}, _T_84};
  assign _T_85 = _GEN_9 << 1;
  assign _T_87 = _T_85 & 32'haaaaaaaa;
  assign _T_88 = _T_83 | _T_87;
  assign shin = _T_37 ? io_in1 : _T_88;
  assign _T_90 = shin[31];
  assign _T_91 = _T_9 & _T_90;
  assign _T_92 = {_T_91,shin};
  assign _T_93 = $signed(_T_92);
  assign _T_94 = $signed(_T_93) >>> shamt;
  assign shout_r = _T_94[31:0];
  assign _T_99 = shout_r[31:16];
  assign _T_100 = {{16'd0}, _T_99};
  assign _T_101 = shout_r[15:0];
  assign _GEN_10 = {{16'd0}, _T_101};
  assign _T_102 = _GEN_10 << 16;
  assign _T_104 = _T_102 & 32'hffff0000;
  assign _T_105 = _T_100 | _T_104;
  assign _T_109 = _T_105[31:8];
  assign _GEN_11 = {{8'd0}, _T_109};
  assign _T_110 = _GEN_11 & 32'hff00ff;
  assign _T_111 = _T_105[23:0];
  assign _GEN_12 = {{8'd0}, _T_111};
  assign _T_112 = _GEN_12 << 8;
  assign _T_114 = _T_112 & 32'hff00ff00;
  assign _T_115 = _T_110 | _T_114;
  assign _T_119 = _T_115[31:4];
  assign _GEN_13 = {{4'd0}, _T_119};
  assign _T_120 = _GEN_13 & 32'hf0f0f0f;
  assign _T_121 = _T_115[27:0];
  assign _GEN_14 = {{4'd0}, _T_121};
  assign _T_122 = _GEN_14 << 4;
  assign _T_124 = _T_122 & 32'hf0f0f0f0;
  assign _T_125 = _T_120 | _T_124;
  assign _T_129 = _T_125[31:2];
  assign _GEN_15 = {{2'd0}, _T_129};
  assign _T_130 = _GEN_15 & 32'h33333333;
  assign _T_131 = _T_125[29:0];
  assign _GEN_16 = {{2'd0}, _T_131};
  assign _T_132 = _GEN_16 << 2;
  assign _T_134 = _T_132 & 32'hcccccccc;
  assign _T_135 = _T_130 | _T_134;
  assign _T_139 = _T_135[31:1];
  assign _GEN_17 = {{1'd0}, _T_139};
  assign _T_140 = _GEN_17 & 32'h55555555;
  assign _T_141 = _T_135[30:0];
  assign _GEN_18 = {{1'd0}, _T_141};
  assign _T_142 = _GEN_18 << 1;
  assign _T_144 = _T_142 & 32'haaaaaaaa;
  assign shout_l = _T_140 | _T_144;
  assign _T_151 = _T_37 ? shout_r : 32'h0;
  assign _T_153 = io_fn == 4'h1;
  assign _T_155 = _T_153 ? shout_l : 32'h0;
  assign shout = _T_151 | _T_155;
  assign _T_157 = io_fn == 4'h4;
  assign _T_159 = io_fn == 4'h6;
  assign _T_160 = _T_157 | _T_159;
  assign _T_162 = _T_160 ? in1_xor_in2 : 32'h0;
  assign _T_166 = io_fn == 4'h7;
  assign _T_167 = _T_159 | _T_166;
  assign _T_168 = io_in1 & io_in2;
  assign _T_170 = _T_167 ? _T_168 : 32'h0;
  assign logic$ = _T_162 | _T_170;
  assign _T_172 = io_fn == 4'h2;
  assign _T_174 = io_fn == 4'h3;
  assign _T_175 = _T_172 | _T_174;
  assign _T_177 = io_fn >= 4'hc;
  assign _T_178 = _T_175 | _T_177;
  assign _T_179 = _T_178 & io_cmp_out;
  assign _GEN_19 = {{31'd0}, _T_179};
  assign _T_180 = _GEN_19 | logic$;
  assign shift_logic = _T_180 | shout;
  assign _T_182 = io_fn == 4'h0;
  assign _T_184 = io_fn == 4'ha;
  assign _T_185 = _T_182 | _T_184;
  assign out = _T_185 ? io_adder_out : shift_logic;
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [3:0]  io_req_bits_fn,
  input  [31:0] io_req_bits_in1,
  input  [31:0] io_req_bits_in2,
  input  [4:0]  io_req_bits_tag,
  input         io_kill,
  input         io_resp_ready,
  output        io_resp_valid,
  output [31:0] io_resp_bits_data,
  output [4:0]  io_resp_bits_tag
);
  reg [2:0] state;
  reg [31:0] _RAND_0;
  reg [4:0] req_tag;
  reg [31:0] _RAND_1;
  reg [5:0] count;
  reg [31:0] _RAND_2;
  reg  neg_out;
  reg [31:0] _RAND_3;
  reg  isHi;
  reg [31:0] _RAND_4;
  reg  resHi;
  reg [31:0] _RAND_5;
  reg [32:0] divisor;
  reg [63:0] _RAND_6;
  reg [65:0] remainder;
  reg [95:0] _RAND_7;
  wire [3:0] _T_32;
  wire  _T_34;
  wire [3:0] _T_36;
  wire  _T_38;
  wire  _T_41;
  wire [3:0] _T_43;
  wire  _T_45;
  wire [3:0] _T_47;
  wire  _T_49;
  wire  _T_52;
  wire  _T_53;
  wire [3:0] _T_55;
  wire  _T_57;
  wire [3:0] _T_59;
  wire  _T_61;
  wire  _T_64;
  wire  _T_65;
  wire  _T_74;
  wire  lhs_sign;
  wire [15:0] _T_80;
  wire [15:0] _T_82;
  wire [31:0] lhs_in;
  wire  _T_88;
  wire  rhs_sign;
  wire [15:0] _T_94;
  wire [15:0] _T_96;
  wire [31:0] rhs_in;
  wire [32:0] _T_97;
  wire [33:0] _T_98;
  wire [33:0] _T_99;
  wire [32:0] subtractor;
  wire [31:0] _T_100;
  wire [31:0] _T_101;
  wire [31:0] result;
  wire [32:0] _T_103;
  wire [32:0] _T_104;
  wire [31:0] negated_remainder;
  wire  _T_105;
  wire  _T_106;
  wire [65:0] _GEN_0;
  wire  _T_107;
  wire [32:0] _GEN_1;
  wire [65:0] _GEN_2;
  wire [32:0] _GEN_3;
  wire [2:0] _GEN_4;
  wire  _T_108;
  wire [65:0] _GEN_5;
  wire [2:0] _GEN_6;
  wire  _GEN_7;
  wire  _T_110;
  wire [32:0] _T_111;
  wire [64:0] _T_113;
  wire  _T_114;
  wire [31:0] _T_115;
  wire [32:0] _T_116;
  wire [32:0] _T_117;
  wire [32:0] _T_118;
  wire [7:0] _T_119;
  wire [8:0] _T_120;
  wire [8:0] _T_121;
  wire [32:0] _GEN_35;
  wire [41:0] _T_122;
  wire [41:0] _GEN_36;
  wire [42:0] _T_123;
  wire [41:0] _T_124;
  wire [41:0] _T_125;
  wire [23:0] _T_126;
  wire [41:0] _T_127;
  wire [65:0] _T_128;
  wire  _T_130;
  wire  _T_131;
  wire  _T_146;
  wire [32:0] _T_161;
  wire [31:0] _T_163;
  wire [64:0] _T_164;
  wire [32:0] _T_165;
  wire [31:0] _T_166;
  wire [33:0] _T_167;
  wire [65:0] _T_168;
  wire [6:0] _T_170;
  wire [5:0] _T_171;
  wire  _T_173;
  wire [2:0] _GEN_8;
  wire  _GEN_9;
  wire [65:0] _GEN_10;
  wire [5:0] _GEN_11;
  wire [2:0] _GEN_12;
  wire  _GEN_13;
  wire  _T_175;
  wire  _T_176;
  wire [31:0] _T_177;
  wire [31:0] _T_178;
  wire [31:0] _T_179;
  wire  _T_182;
  wire [63:0] _T_183;
  wire [64:0] _T_184;
  wire  _T_186;
  wire [2:0] _T_187;
  wire [2:0] _GEN_14;
  wire  _GEN_15;
  wire  _T_192;
  wire  _T_196;
  wire  _T_199;
  wire  _GEN_16;
  wire [65:0] _GEN_17;
  wire [2:0] _GEN_18;
  wire  _GEN_19;
  wire [5:0] _GEN_20;
  wire  _GEN_21;
  wire  _T_201;
  wire  _T_202;
  wire [2:0] _GEN_22;
  wire  _T_203;
  wire  _T_204;
  wire [2:0] _T_205;
  wire [2:0] _T_206;
  wire  _T_218;
  wire  _T_219;
  wire [32:0] _T_220;
  wire [2:0] _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire [5:0] _GEN_26;
  wire  _GEN_27;
  wire [32:0] _GEN_28;
  wire [65:0] _GEN_29;
  wire [4:0] _GEN_34;
  wire [15:0] _T_232;
  wire [15:0] _T_233;
  wire [31:0] _T_244;
  wire  _T_245;
  wire  _T_246;
  wire  _T_247;
  wire  _T_248;
  assign io_req_ready = _T_248;
  assign io_resp_valid = _T_247;
  assign io_resp_bits_data = _T_244;
  assign io_resp_bits_tag = req_tag;
  assign _T_32 = io_req_bits_fn & 4'h4;
  assign _T_34 = _T_32 == 4'h0;
  assign _T_36 = io_req_bits_fn & 4'h8;
  assign _T_38 = _T_36 == 4'h8;
  assign _T_41 = _T_34 | _T_38;
  assign _T_43 = io_req_bits_fn & 4'h5;
  assign _T_45 = _T_43 == 4'h1;
  assign _T_47 = io_req_bits_fn & 4'h2;
  assign _T_49 = _T_47 == 4'h2;
  assign _T_52 = _T_45 | _T_49;
  assign _T_53 = _T_52 | _T_38;
  assign _T_55 = io_req_bits_fn & 4'h9;
  assign _T_57 = _T_55 == 4'h0;
  assign _T_59 = io_req_bits_fn & 4'h3;
  assign _T_61 = _T_59 == 4'h0;
  assign _T_64 = _T_57 | _T_34;
  assign _T_65 = _T_64 | _T_61;
  assign _T_74 = io_req_bits_in1[31];
  assign lhs_sign = _T_65 & _T_74;
  assign _T_80 = io_req_bits_in1[31:16];
  assign _T_82 = io_req_bits_in1[15:0];
  assign lhs_in = {_T_80,_T_82};
  assign _T_88 = io_req_bits_in2[31];
  assign rhs_sign = _T_64 & _T_88;
  assign _T_94 = io_req_bits_in2[31:16];
  assign _T_96 = io_req_bits_in2[15:0];
  assign rhs_in = {_T_94,_T_96};
  assign _T_97 = remainder[64:32];
  assign _T_98 = _T_97 - divisor;
  assign _T_99 = $unsigned(_T_98);
  assign subtractor = _T_99[32:0];
  assign _T_100 = remainder[64:33];
  assign _T_101 = remainder[31:0];
  assign result = resHi ? _T_100 : _T_101;
  assign _T_103 = 32'h0 - result;
  assign _T_104 = $unsigned(_T_103);
  assign negated_remainder = _T_104[31:0];
  assign _T_105 = state == 3'h1;
  assign _T_106 = remainder[31];
  assign _GEN_0 = _T_106 ? {{34'd0}, negated_remainder} : remainder;
  assign _T_107 = divisor[31];
  assign _GEN_1 = _T_107 ? subtractor : divisor;
  assign _GEN_2 = _T_105 ? _GEN_0 : remainder;
  assign _GEN_3 = _T_105 ? _GEN_1 : divisor;
  assign _GEN_4 = _T_105 ? 3'h3 : state;
  assign _T_108 = state == 3'h5;
  assign _GEN_5 = _T_108 ? {{34'd0}, negated_remainder} : _GEN_2;
  assign _GEN_6 = _T_108 ? 3'h7 : _GEN_4;
  assign _GEN_7 = _T_108 ? 1'h0 : resHi;
  assign _T_110 = state == 3'h2;
  assign _T_111 = remainder[65:33];
  assign _T_113 = {_T_111,_T_101};
  assign _T_114 = remainder[32];
  assign _T_115 = _T_113[31:0];
  assign _T_116 = _T_113[64:32];
  assign _T_117 = $signed(_T_116);
  assign _T_118 = $signed(divisor);
  assign _T_119 = _T_115[7:0];
  assign _T_120 = {_T_114,_T_119};
  assign _T_121 = $signed(_T_120);
  assign _GEN_35 = {{24{_T_121[8]}},_T_121};
  assign _T_122 = $signed(_GEN_35) * $signed(_T_118);
  assign _GEN_36 = {{9{_T_117[32]}},_T_117};
  assign _T_123 = $signed(_T_122) + $signed(_GEN_36);
  assign _T_124 = _T_123[41:0];
  assign _T_125 = $signed(_T_124);
  assign _T_126 = _T_115[31:8];
  assign _T_127 = $unsigned(_T_125);
  assign _T_128 = {_T_127,_T_126};
  assign _T_130 = count == 6'h2;
  assign _T_131 = _T_130 & neg_out;
  assign _T_146 = isHi == 1'h0;
  assign _T_161 = _T_128[64:32];
  assign _T_163 = _T_128[31:0];
  assign _T_164 = {_T_161,_T_163};
  assign _T_165 = _T_164[64:32];
  assign _T_166 = _T_164[31:0];
  assign _T_167 = {_T_165,_T_131};
  assign _T_168 = {_T_167,_T_166};
  assign _T_170 = count + 6'h1;
  assign _T_171 = _T_170[5:0];
  assign _T_173 = count == 6'h3;
  assign _GEN_8 = _T_173 ? 3'h6 : _GEN_6;
  assign _GEN_9 = _T_173 ? isHi : _GEN_7;
  assign _GEN_10 = _T_110 ? _T_168 : _GEN_5;
  assign _GEN_11 = _T_110 ? _T_171 : count;
  assign _GEN_12 = _T_110 ? _GEN_8 : _GEN_6;
  assign _GEN_13 = _T_110 ? _GEN_9 : _GEN_7;
  assign _T_175 = state == 3'h3;
  assign _T_176 = subtractor[32];
  assign _T_177 = remainder[63:32];
  assign _T_178 = subtractor[31:0];
  assign _T_179 = _T_176 ? _T_177 : _T_178;
  assign _T_182 = _T_176 == 1'h0;
  assign _T_183 = {_T_179,_T_101};
  assign _T_184 = {_T_183,_T_182};
  assign _T_186 = count == 6'h20;
  assign _T_187 = neg_out ? 3'h5 : 3'h7;
  assign _GEN_14 = _T_186 ? _T_187 : _GEN_12;
  assign _GEN_15 = _T_186 ? isHi : _GEN_13;
  assign _T_192 = count == 6'h0;
  assign _T_196 = _T_192 & _T_182;
  assign _T_199 = _T_196 & _T_146;
  assign _GEN_16 = _T_199 ? 1'h0 : neg_out;
  assign _GEN_17 = _T_175 ? {{1'd0}, _T_184} : _GEN_10;
  assign _GEN_18 = _T_175 ? _GEN_14 : _GEN_12;
  assign _GEN_19 = _T_175 ? _GEN_15 : _GEN_13;
  assign _GEN_20 = _T_175 ? _T_171 : _GEN_11;
  assign _GEN_21 = _T_175 ? _GEN_16 : neg_out;
  assign _T_201 = io_resp_ready & io_resp_valid;
  assign _T_202 = _T_201 | io_kill;
  assign _GEN_22 = _T_202 ? 3'h0 : _GEN_18;
  assign _T_203 = io_req_ready & io_req_valid;
  assign _T_204 = lhs_sign | rhs_sign;
  assign _T_205 = _T_204 ? 3'h1 : 3'h3;
  assign _T_206 = _T_41 ? 3'h2 : _T_205;
  assign _T_218 = lhs_sign != rhs_sign;
  assign _T_219 = _T_53 ? lhs_sign : _T_218;
  assign _T_220 = {rhs_sign,rhs_in};
  assign _GEN_23 = _T_203 ? _T_206 : _GEN_22;
  assign _GEN_24 = _T_203 ? _T_53 : isHi;
  assign _GEN_25 = _T_203 ? 1'h0 : _GEN_19;
  assign _GEN_26 = _T_203 ? 6'h0 : _GEN_20;
  assign _GEN_27 = _T_203 ? _T_219 : _GEN_21;
  assign _GEN_28 = _T_203 ? _T_220 : _GEN_3;
  assign _GEN_29 = _T_203 ? {{34'd0}, lhs_in} : _GEN_17;
  assign _GEN_34 = _T_203 ? io_req_bits_tag : req_tag;
  assign _T_232 = result[31:16];
  assign _T_233 = result[15:0];
  assign _T_244 = {_T_232,_T_233};
  assign _T_245 = state == 3'h6;
  assign _T_246 = state == 3'h7;
  assign _T_247 = _T_245 | _T_246;
  assign _T_248 = state == 3'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  req_tag = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  count = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  neg_out = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  isHi = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  resHi = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{$random}};
  divisor = _RAND_6[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{$random}};
  remainder = _RAND_7[65:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_203) begin
        if (_T_41) begin
          state <= 3'h2;
        end else begin
          if (_T_204) begin
            state <= 3'h1;
          end else begin
            state <= 3'h3;
          end
        end
      end else begin
        if (_T_202) begin
          state <= 3'h0;
        end else begin
          if (_T_175) begin
            if (_T_186) begin
              if (neg_out) begin
                state <= 3'h5;
              end else begin
                state <= 3'h7;
              end
            end else begin
              if (_T_110) begin
                if (_T_173) begin
                  state <= 3'h6;
                end else begin
                  if (_T_108) begin
                    state <= 3'h7;
                  end else begin
                    if (_T_105) begin
                      state <= 3'h3;
                    end
                  end
                end
              end else begin
                if (_T_108) begin
                  state <= 3'h7;
                end else begin
                  if (_T_105) begin
                    state <= 3'h3;
                  end
                end
              end
            end
          end else begin
            if (_T_110) begin
              if (_T_173) begin
                state <= 3'h6;
              end else begin
                if (_T_108) begin
                  state <= 3'h7;
                end else begin
                  if (_T_105) begin
                    state <= 3'h3;
                  end
                end
              end
            end else begin
              if (_T_108) begin
                state <= 3'h7;
              end else begin
                if (_T_105) begin
                  state <= 3'h3;
                end
              end
            end
          end
        end
      end
    end
    if (_T_203) begin
      req_tag <= io_req_bits_tag;
    end
    if (_T_203) begin
      count <= 6'h0;
    end else begin
      if (_T_175) begin
        count <= _T_171;
      end else begin
        if (_T_110) begin
          count <= _T_171;
        end
      end
    end
    if (_T_203) begin
      if (_T_53) begin
        neg_out <= lhs_sign;
      end else begin
        neg_out <= _T_218;
      end
    end else begin
      if (_T_175) begin
        if (_T_199) begin
          neg_out <= 1'h0;
        end
      end
    end
    if (_T_203) begin
      isHi <= _T_53;
    end
    if (_T_203) begin
      resHi <= 1'h0;
    end else begin
      if (_T_175) begin
        if (_T_186) begin
          resHi <= isHi;
        end else begin
          if (_T_110) begin
            if (_T_173) begin
              resHi <= isHi;
            end else begin
              if (_T_108) begin
                resHi <= 1'h0;
              end
            end
          end else begin
            if (_T_108) begin
              resHi <= 1'h0;
            end
          end
        end
      end else begin
        if (_T_110) begin
          if (_T_173) begin
            resHi <= isHi;
          end else begin
            if (_T_108) begin
              resHi <= 1'h0;
            end
          end
        end else begin
          if (_T_108) begin
            resHi <= 1'h0;
          end
        end
      end
    end
    if (_T_203) begin
      divisor <= _T_220;
    end else begin
      if (_T_105) begin
        if (_T_107) begin
          divisor <= subtractor;
        end
      end
    end
    if (_T_203) begin
      remainder <= {{34'd0}, lhs_in};
    end else begin
      if (_T_175) begin
        remainder <= {{1'd0}, _T_184};
      end else begin
        if (_T_110) begin
          remainder <= _T_168;
        end else begin
          if (_T_108) begin
            remainder <= {{34'd0}, negated_remainder};
          end else begin
            if (_T_105) begin
              if (_T_106) begin
                remainder <= {{34'd0}, negated_remainder};
              end
            end
          end
        end
      end
    end
  end
endmodule
module Rocket(
  input         clock,
  input         reset,
  input         io_hartid,
  input         io_interrupts_debug,
  input         io_interrupts_mtip,
  input         io_interrupts_msip,
  input         io_interrupts_meip,
  output        io_imem_req_valid,
  output [31:0] io_imem_req_bits_pc,
  output        io_imem_req_bits_speculative,
  output        io_imem_sfence_valid,
  output        io_imem_sfence_bits_rs1,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input         io_imem_resp_bits_btb_valid,
  input         io_imem_resp_bits_btb_bits_taken,
  input         io_imem_resp_bits_btb_bits_bridx,
  input  [31:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data,
  input         io_imem_resp_bits_xcpt_pf_inst,
  input         io_imem_resp_bits_xcpt_ae_inst,
  input         io_imem_resp_bits_replay,
  output        io_imem_flush_icache,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [6:0]  io_dmem_req_bits_tag,
  output [4:0]  io_dmem_req_bits_cmd,
  output [2:0]  io_dmem_req_bits_typ,
  output        io_dmem_req_bits_phys,
  output        io_dmem_s1_kill,
  output [31:0] io_dmem_s1_data_data,
  output [3:0]  io_dmem_s1_data_mask,
  input         io_dmem_s2_nack,
  input         io_dmem_resp_valid,
  input  [6:0]  io_dmem_resp_bits_tag,
  input  [31:0] io_dmem_resp_bits_data,
  input         io_dmem_resp_bits_replay,
  input         io_dmem_resp_bits_has_data,
  input  [31:0] io_dmem_resp_bits_data_word_bypass,
  input         io_dmem_replay_next,
  input         io_dmem_s2_xcpt_ma_ld,
  input         io_dmem_s2_xcpt_ma_st,
  input         io_dmem_s2_xcpt_pf_ld,
  input         io_dmem_s2_xcpt_pf_st,
  input         io_dmem_s2_xcpt_ae_ld,
  input         io_dmem_s2_xcpt_ae_st,
  output        io_dmem_invalidate_lr,
  input         io_dmem_ordered,
  output [21:0] io_ptw_ptbr_ppn,
  output        io_ptw_sfence_valid,
  output        io_ptw_sfence_bits_rs1,
  output [1:0]  io_ptw_status_dprv,
  output [1:0]  io_ptw_status_prv,
  output        io_ptw_status_mxr,
  output        io_ptw_status_sum,
  output        io_ptw_pmp_0_cfg_l,
  output [1:0]  io_ptw_pmp_0_cfg_a,
  output        io_ptw_pmp_0_cfg_x,
  output        io_ptw_pmp_0_cfg_w,
  output        io_ptw_pmp_0_cfg_r,
  output [29:0] io_ptw_pmp_0_addr,
  output [31:0] io_ptw_pmp_0_mask,
  output        io_ptw_pmp_1_cfg_l,
  output [1:0]  io_ptw_pmp_1_cfg_a,
  output        io_ptw_pmp_1_cfg_x,
  output        io_ptw_pmp_1_cfg_w,
  output        io_ptw_pmp_1_cfg_r,
  output [29:0] io_ptw_pmp_1_addr,
  output [31:0] io_ptw_pmp_1_mask,
  output        io_ptw_pmp_2_cfg_l,
  output [1:0]  io_ptw_pmp_2_cfg_a,
  output        io_ptw_pmp_2_cfg_x,
  output        io_ptw_pmp_2_cfg_w,
  output        io_ptw_pmp_2_cfg_r,
  output [29:0] io_ptw_pmp_2_addr,
  output [31:0] io_ptw_pmp_2_mask,
  output        io_ptw_pmp_3_cfg_l,
  output [1:0]  io_ptw_pmp_3_cfg_a,
  output        io_ptw_pmp_3_cfg_x,
  output        io_ptw_pmp_3_cfg_w,
  output        io_ptw_pmp_3_cfg_r,
  output [29:0] io_ptw_pmp_3_addr,
  output [31:0] io_ptw_pmp_3_mask,
  output        io_ptw_pmp_4_cfg_l,
  output [1:0]  io_ptw_pmp_4_cfg_a,
  output        io_ptw_pmp_4_cfg_x,
  output        io_ptw_pmp_4_cfg_w,
  output        io_ptw_pmp_4_cfg_r,
  output [29:0] io_ptw_pmp_4_addr,
  output [31:0] io_ptw_pmp_4_mask,
  output        io_ptw_pmp_5_cfg_l,
  output [1:0]  io_ptw_pmp_5_cfg_a,
  output        io_ptw_pmp_5_cfg_x,
  output        io_ptw_pmp_5_cfg_w,
  output        io_ptw_pmp_5_cfg_r,
  output [29:0] io_ptw_pmp_5_addr,
  output [31:0] io_ptw_pmp_5_mask,
  output        io_ptw_pmp_6_cfg_l,
  output [1:0]  io_ptw_pmp_6_cfg_a,
  output        io_ptw_pmp_6_cfg_x,
  output        io_ptw_pmp_6_cfg_w,
  output        io_ptw_pmp_6_cfg_r,
  output [29:0] io_ptw_pmp_6_addr,
  output [31:0] io_ptw_pmp_6_mask,
  output        io_ptw_pmp_7_cfg_l,
  output [1:0]  io_ptw_pmp_7_cfg_a,
  output        io_ptw_pmp_7_cfg_x,
  output        io_ptw_pmp_7_cfg_w,
  output        io_ptw_pmp_7_cfg_r,
  output [29:0] io_ptw_pmp_7_addr,
  output [31:0] io_ptw_pmp_7_mask,
  input  [31:0] io_fpu_store_data,
  input  [31:0] io_fpu_toint_data,
  input         io_fpu_nack_mem,
  input         io_fpu_dec_wen,
  input         io_fpu_dec_ren1,
  input         io_fpu_dec_ren2,
  input         io_fpu_dec_ren3,
  input         io_rocc_cmd_ready,
  input         io_rocc_interrupt
);
  reg  ex_ctrl_fp;
  reg [31:0] _RAND_0;
  reg  ex_ctrl_rocc;
  reg [31:0] _RAND_1;
  reg  ex_ctrl_branch;
  reg [31:0] _RAND_2;
  reg  ex_ctrl_jal;
  reg [31:0] _RAND_3;
  reg  ex_ctrl_jalr;
  reg [31:0] _RAND_4;
  reg  ex_ctrl_rxs2;
  reg [31:0] _RAND_5;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [31:0] _RAND_6;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [31:0] _RAND_7;
  reg [2:0] ex_ctrl_sel_imm;
  reg [31:0] _RAND_8;
  reg [3:0] ex_ctrl_alu_fn;
  reg [31:0] _RAND_9;
  reg  ex_ctrl_mem;
  reg [31:0] _RAND_10;
  reg [4:0] ex_ctrl_mem_cmd;
  reg [31:0] _RAND_11;
  reg [2:0] ex_ctrl_mem_type;
  reg [31:0] _RAND_12;
  reg  ex_ctrl_wfd;
  reg [31:0] _RAND_13;
  reg  ex_ctrl_div;
  reg [31:0] _RAND_14;
  reg  ex_ctrl_wxd;
  reg [31:0] _RAND_15;
  reg [2:0] ex_ctrl_csr;
  reg [31:0] _RAND_16;
  reg  ex_ctrl_fence_i;
  reg [31:0] _RAND_17;
  reg  mem_ctrl_fp;
  reg [31:0] _RAND_18;
  reg  mem_ctrl_rocc;
  reg [31:0] _RAND_19;
  reg  mem_ctrl_branch;
  reg [31:0] _RAND_20;
  reg  mem_ctrl_jal;
  reg [31:0] _RAND_21;
  reg  mem_ctrl_jalr;
  reg [31:0] _RAND_22;
  reg  mem_ctrl_mem;
  reg [31:0] _RAND_23;
  reg [2:0] mem_ctrl_mem_type;
  reg [31:0] _RAND_24;
  reg  mem_ctrl_wfd;
  reg [31:0] _RAND_25;
  reg  mem_ctrl_div;
  reg [31:0] _RAND_26;
  reg  mem_ctrl_wxd;
  reg [31:0] _RAND_27;
  reg [2:0] mem_ctrl_csr;
  reg [31:0] _RAND_28;
  reg  mem_ctrl_fence_i;
  reg [31:0] _RAND_29;
  reg  wb_ctrl_rocc;
  reg [31:0] _RAND_30;
  reg  wb_ctrl_mem;
  reg [31:0] _RAND_31;
  reg [2:0] wb_ctrl_mem_type;
  reg [31:0] _RAND_32;
  reg  wb_ctrl_wfd;
  reg [31:0] _RAND_33;
  reg  wb_ctrl_div;
  reg [31:0] _RAND_34;
  reg  wb_ctrl_wxd;
  reg [31:0] _RAND_35;
  reg [2:0] wb_ctrl_csr;
  reg [31:0] _RAND_36;
  reg  wb_ctrl_fence_i;
  reg [31:0] _RAND_37;
  reg  ex_reg_xcpt_interrupt;
  reg [31:0] _RAND_38;
  reg  ex_reg_valid;
  reg [31:0] _RAND_39;
  reg  ex_reg_rvc;
  reg [31:0] _RAND_40;
  reg  ex_reg_xcpt;
  reg [31:0] _RAND_41;
  reg  ex_reg_flush_pipe;
  reg [31:0] _RAND_42;
  reg  ex_reg_load_use;
  reg [31:0] _RAND_43;
  reg [31:0] ex_cause;
  reg [31:0] _RAND_44;
  reg  ex_reg_replay;
  reg [31:0] _RAND_45;
  reg [31:0] ex_reg_pc;
  reg [31:0] _RAND_46;
  reg [31:0] ex_reg_inst;
  reg [31:0] _RAND_47;
  reg  mem_reg_xcpt_interrupt;
  reg [31:0] _RAND_48;
  reg  mem_reg_valid;
  reg [31:0] _RAND_49;
  reg  mem_reg_rvc;
  reg [31:0] _RAND_50;
  reg  mem_reg_xcpt;
  reg [31:0] _RAND_51;
  reg  mem_reg_replay;
  reg [31:0] _RAND_52;
  reg  mem_reg_flush_pipe;
  reg [31:0] _RAND_53;
  reg [31:0] mem_reg_cause;
  reg [31:0] _RAND_54;
  reg  mem_reg_slow_bypass;
  reg [31:0] _RAND_55;
  reg  mem_reg_load;
  reg [31:0] _RAND_56;
  reg  mem_reg_store;
  reg [31:0] _RAND_57;
  reg  mem_reg_sfence;
  reg [31:0] _RAND_58;
  reg [31:0] mem_reg_pc;
  reg [31:0] _RAND_59;
  reg [31:0] mem_reg_inst;
  reg [31:0] _RAND_60;
  reg [31:0] bypass_mux_1;
  reg [31:0] _RAND_61;
  reg [31:0] mem_reg_rs2;
  reg [31:0] _RAND_62;
  reg  wb_reg_valid;
  reg [31:0] _RAND_63;
  reg  wb_reg_rvc;
  reg [31:0] _RAND_64;
  reg  wb_reg_xcpt;
  reg [31:0] _RAND_65;
  reg  wb_reg_replay;
  reg [31:0] _RAND_66;
  reg  wb_reg_flush_pipe;
  reg [31:0] _RAND_67;
  reg [31:0] wb_reg_cause;
  reg [31:0] _RAND_68;
  reg  wb_reg_sfence;
  reg [31:0] _RAND_69;
  reg [31:0] wb_reg_pc;
  reg [31:0] _RAND_70;
  reg [31:0] wb_reg_inst;
  reg [31:0] _RAND_71;
  reg [31:0] bypass_mux_2;
  reg [31:0] _RAND_72;
  wire  take_pc;
  wire  ibuf_clock;
  wire  ibuf_reset;
  wire  ibuf_io_imem_ready;
  wire  ibuf_io_imem_valid;
  wire  ibuf_io_imem_bits_btb_valid;
  wire  ibuf_io_imem_bits_btb_bits_taken;
  wire  ibuf_io_imem_bits_btb_bits_bridx;
  wire [31:0] ibuf_io_imem_bits_pc;
  wire [31:0] ibuf_io_imem_bits_data;
  wire  ibuf_io_imem_bits_xcpt_pf_inst;
  wire  ibuf_io_imem_bits_xcpt_ae_inst;
  wire  ibuf_io_imem_bits_replay;
  wire  ibuf_io_kill;
  wire [31:0] ibuf_io_pc;
  wire  ibuf_io_inst_0_ready;
  wire  ibuf_io_inst_0_valid;
  wire  ibuf_io_inst_0_bits_xcpt0_pf_inst;
  wire  ibuf_io_inst_0_bits_xcpt0_ae_inst;
  wire  ibuf_io_inst_0_bits_xcpt1_pf_inst;
  wire  ibuf_io_inst_0_bits_xcpt1_ae_inst;
  wire  ibuf_io_inst_0_bits_replay;
  wire  ibuf_io_inst_0_bits_rvc;
  wire [31:0] ibuf_io_inst_0_bits_inst_bits;
  wire [4:0] ibuf_io_inst_0_bits_inst_rd;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs1;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs2;
  wire [4:0] ibuf_io_inst_0_bits_inst_rs3;
  wire [31:0] ibuf_io_inst_0_bits_raw;
  wire [31:0] _T_679;
  wire  _T_681;
  wire [31:0] _T_683;
  wire  _T_685;
  wire [31:0] _T_687;
  wire  _T_689;
  wire [31:0] _T_691;
  wire  _T_693;
  wire [31:0] _T_695;
  wire  _T_697;
  wire [31:0] _T_699;
  wire  _T_701;
  wire [31:0] _T_703;
  wire  _T_705;
  wire [31:0] _T_707;
  wire  _T_709;
  wire [31:0] _T_711;
  wire  _T_713;
  wire [31:0] _T_715;
  wire  _T_717;
  wire  _T_721;
  wire [31:0] _T_723;
  wire  _T_725;
  wire  _T_729;
  wire [31:0] _T_731;
  wire  _T_733;
  wire  _T_737;
  wire [31:0] _T_739;
  wire  _T_741;
  wire [31:0] _T_743;
  wire  _T_745;
  wire  _T_747;
  wire  _T_749;
  wire  _T_751;
  wire [31:0] _T_753;
  wire  _T_755;
  wire [31:0] _T_757;
  wire  _T_759;
  wire [31:0] _T_761;
  wire  _T_763;
  wire  _T_767;
  wire  _T_770;
  wire  _T_771;
  wire  _T_772;
  wire  _T_773;
  wire  _T_774;
  wire  _T_775;
  wire  _T_776;
  wire  _T_777;
  wire  _T_778;
  wire  _T_779;
  wire  _T_780;
  wire  _T_781;
  wire  _T_782;
  wire  _T_783;
  wire  _T_784;
  wire  _T_785;
  wire  _T_786;
  wire  _T_787;
  wire  _T_788;
  wire  _T_789;
  wire  _T_790;
  wire  _T_791;
  wire  _T_792;
  wire [31:0] _T_796;
  wire  _T_798;
  wire [31:0] _T_802;
  wire  _T_804;
  wire [31:0] _T_808;
  wire  _T_810;
  wire [31:0] _T_814;
  wire  _T_816;
  wire [31:0] _T_818;
  wire  _T_820;
  wire [31:0] _T_822;
  wire  _T_824;
  wire  _T_827;
  wire  _T_828;
  wire [31:0] _T_830;
  wire  _T_832;
  wire [31:0] _T_834;
  wire  _T_836;
  wire [31:0] _T_838;
  wire  _T_840;
  wire [31:0] _T_842;
  wire  _T_844;
  wire  _T_847;
  wire  _T_848;
  wire  _T_849;
  wire [31:0] _T_851;
  wire  _T_853;
  wire [31:0] _T_855;
  wire  _T_857;
  wire [31:0] _T_859;
  wire  _T_861;
  wire [31:0] _T_863;
  wire  _T_865;
  wire  _T_868;
  wire  _T_869;
  wire  _T_870;
  wire  _T_871;
  wire  _T_875;
  wire [31:0] _T_877;
  wire  _T_879;
  wire  _T_882;
  wire  _T_883;
  wire [1:0] _T_884;
  wire [31:0] _T_886;
  wire  _T_888;
  wire  _T_891;
  wire  _T_892;
  wire  _T_893;
  wire [31:0] _T_895;
  wire  _T_897;
  wire  _T_900;
  wire [1:0] _T_901;
  wire [31:0] _T_903;
  wire  _T_905;
  wire  _T_909;
  wire  _T_912;
  wire  _T_916;
  wire  _T_919;
  wire  _T_923;
  wire [31:0] _T_925;
  wire  _T_927;
  wire  _T_930;
  wire  _T_931;
  wire [1:0] _T_932;
  wire [2:0] _T_933;
  wire [31:0] _T_941;
  wire  _T_943;
  wire [31:0] _T_945;
  wire  _T_947;
  wire [31:0] _T_949;
  wire  _T_951;
  wire  _T_954;
  wire  _T_955;
  wire [31:0] _T_957;
  wire  _T_959;
  wire [31:0] _T_961;
  wire  _T_963;
  wire [31:0] _T_965;
  wire  _T_967;
  wire [31:0] _T_969;
  wire  _T_971;
  wire [31:0] _T_973;
  wire  _T_975;
  wire [31:0] _T_977;
  wire  _T_979;
  wire  _T_982;
  wire  _T_983;
  wire  _T_984;
  wire  _T_985;
  wire  _T_986;
  wire [31:0] _T_988;
  wire  _T_990;
  wire [31:0] _T_992;
  wire  _T_994;
  wire [31:0] _T_996;
  wire  _T_998;
  wire [31:0] _T_1000;
  wire  _T_1002;
  wire  _T_1005;
  wire  _T_1006;
  wire  _T_1007;
  wire [31:0] _T_1009;
  wire  _T_1011;
  wire [31:0] _T_1013;
  wire  _T_1015;
  wire  _T_1018;
  wire  _T_1019;
  wire  _T_1020;
  wire [1:0] _T_1021;
  wire [1:0] _T_1022;
  wire [3:0] _T_1023;
  wire [31:0] _T_1025;
  wire  _T_1027;
  wire [31:0] _T_1029;
  wire  _T_1031;
  wire  _T_1034;
  wire  _T_1035;
  wire  _T_1036;
  wire  _T_1037;
  wire  _T_1038;
  wire  _T_1039;
  wire [31:0] _T_1041;
  wire  _T_1043;
  wire [31:0] _T_1045;
  wire  _T_1047;
  wire [31:0] _T_1049;
  wire  _T_1051;
  wire [31:0] _T_1053;
  wire  _T_1055;
  wire  _T_1058;
  wire  _T_1059;
  wire  _T_1060;
  wire [31:0] _T_1062;
  wire  _T_1064;
  wire [31:0] _T_1066;
  wire  _T_1068;
  wire  _T_1071;
  wire [31:0] _T_1073;
  wire  _T_1075;
  wire [31:0] _T_1077;
  wire  _T_1079;
  wire [31:0] _T_1081;
  wire  _T_1083;
  wire  _T_1086;
  wire  _T_1087;
  wire  _T_1088;
  wire [31:0] _T_1090;
  wire  _T_1092;
  wire [1:0] _T_1096;
  wire [1:0] _T_1097;
  wire [2:0] _T_1098;
  wire [4:0] _T_1099;
  wire [31:0] _T_1101;
  wire  _T_1103;
  wire [31:0] _T_1107;
  wire  _T_1109;
  wire [31:0] _T_1113;
  wire  _T_1115;
  wire [1:0] _T_1118;
  wire [2:0] _T_1119;
  wire [31:0] _T_1125;
  wire  _T_1127;
  wire  _T_1133;
  wire  _T_1137;
  wire [31:0] _T_1139;
  wire  _T_1141;
  wire  _T_1145;
  wire [31:0] _T_1147;
  wire  _T_1149;
  wire  _T_1152;
  wire  _T_1153;
  wire  _T_1154;
  wire  _T_1155;
  wire  _T_1156;
  wire  _T_1157;
  wire [31:0] _T_1159;
  wire  _T_1161;
  wire  _T_1167;
  wire [31:0] _T_1171;
  wire  _T_1173;
  wire [1:0] _T_1176;
  wire [2:0] _T_1177;
  wire [31:0] _T_1179;
  wire  _T_1181;
  wire [31:0] _T_1185;
  wire  _T_1187;
  wire [31:0] _T_1191;
  wire  _T_1193;
  reg  id_reg_fence;
  reg [31:0] _RAND_73;
  reg [31:0] _T_1202 [0:30];
  reg [31:0] _RAND_74;
  wire [31:0] _T_1202__T_1211_data;
  wire [4:0] _T_1202__T_1211_addr;
  reg [31:0] _RAND_75;
  wire [31:0] _T_1202__T_1221_data;
  wire [4:0] _T_1202__T_1221_addr;
  reg [31:0] _RAND_76;
  wire [31:0] _T_1202__T_2124_data;
  wire [4:0] _T_1202__T_2124_addr;
  wire  _T_1202__T_2124_mask;
  wire  _T_1202__T_2124_en;
  wire  _T_1206;
  wire [4:0] _T_1209;
  wire [4:0] _T_1210;
  wire [31:0] _T_1212;
  wire [4:0] _T_1219;
  wire [4:0] _T_1220;
  wire [31:0] _T_1222;
  wire  csr_clock;
  wire  csr_reset;
  wire  csr_io_interrupts_debug;
  wire  csr_io_interrupts_mtip;
  wire  csr_io_interrupts_msip;
  wire  csr_io_interrupts_meip;
  wire  csr_io_hartid;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [31:0] csr_io_rw_rdata;
  wire [31:0] csr_io_rw_wdata;
  wire [11:0] csr_io_decode_csr;
  wire  csr_io_decode_read_illegal;
  wire  csr_io_decode_write_illegal;
  wire  csr_io_decode_write_flush;
  wire  csr_io_decode_system_illegal;
  wire  csr_io_csr_stall;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire [31:0] csr_io_status_isa;
  wire [1:0] csr_io_status_dprv;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [26:0] csr_io_status_zero2;
  wire [1:0] csr_io_status_sxl;
  wire [1:0] csr_io_status_uxl;
  wire  csr_io_status_sd_rv32;
  wire [7:0] csr_io_status_zero1;
  wire  csr_io_status_tsr;
  wire  csr_io_status_tw;
  wire  csr_io_status_tvm;
  wire  csr_io_status_mxr;
  wire  csr_io_status_sum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [21:0] csr_io_ptbr_ppn;
  wire [31:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire [31:0] csr_io_cause;
  wire [31:0] csr_io_pc;
  wire [31:0] csr_io_badaddr;
  wire [31:0] csr_io_time;
  wire  csr_io_rocc_interrupt;
  wire  csr_io_interrupt;
  wire [31:0] csr_io_interrupt_cause;
  wire  csr_io_bp_0_control_action;
  wire  csr_io_bp_0_control_chain;
  wire [1:0] csr_io_bp_0_control_tmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_h;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_x;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_r;
  wire [31:0] csr_io_bp_0_address;
  wire  csr_io_pmp_0_cfg_l;
  wire [1:0] csr_io_pmp_0_cfg_a;
  wire  csr_io_pmp_0_cfg_x;
  wire  csr_io_pmp_0_cfg_w;
  wire  csr_io_pmp_0_cfg_r;
  wire [29:0] csr_io_pmp_0_addr;
  wire [31:0] csr_io_pmp_0_mask;
  wire  csr_io_pmp_1_cfg_l;
  wire [1:0] csr_io_pmp_1_cfg_a;
  wire  csr_io_pmp_1_cfg_x;
  wire  csr_io_pmp_1_cfg_w;
  wire  csr_io_pmp_1_cfg_r;
  wire [29:0] csr_io_pmp_1_addr;
  wire [31:0] csr_io_pmp_1_mask;
  wire  csr_io_pmp_2_cfg_l;
  wire [1:0] csr_io_pmp_2_cfg_a;
  wire  csr_io_pmp_2_cfg_x;
  wire  csr_io_pmp_2_cfg_w;
  wire  csr_io_pmp_2_cfg_r;
  wire [29:0] csr_io_pmp_2_addr;
  wire [31:0] csr_io_pmp_2_mask;
  wire  csr_io_pmp_3_cfg_l;
  wire [1:0] csr_io_pmp_3_cfg_a;
  wire  csr_io_pmp_3_cfg_x;
  wire  csr_io_pmp_3_cfg_w;
  wire  csr_io_pmp_3_cfg_r;
  wire [29:0] csr_io_pmp_3_addr;
  wire [31:0] csr_io_pmp_3_mask;
  wire  csr_io_pmp_4_cfg_l;
  wire [1:0] csr_io_pmp_4_cfg_a;
  wire  csr_io_pmp_4_cfg_x;
  wire  csr_io_pmp_4_cfg_w;
  wire  csr_io_pmp_4_cfg_r;
  wire [29:0] csr_io_pmp_4_addr;
  wire [31:0] csr_io_pmp_4_mask;
  wire  csr_io_pmp_5_cfg_l;
  wire [1:0] csr_io_pmp_5_cfg_a;
  wire  csr_io_pmp_5_cfg_x;
  wire  csr_io_pmp_5_cfg_w;
  wire  csr_io_pmp_5_cfg_r;
  wire [29:0] csr_io_pmp_5_addr;
  wire [31:0] csr_io_pmp_5_mask;
  wire  csr_io_pmp_6_cfg_l;
  wire [1:0] csr_io_pmp_6_cfg_a;
  wire  csr_io_pmp_6_cfg_x;
  wire  csr_io_pmp_6_cfg_w;
  wire  csr_io_pmp_6_cfg_r;
  wire [29:0] csr_io_pmp_6_addr;
  wire [31:0] csr_io_pmp_6_mask;
  wire  csr_io_pmp_7_cfg_l;
  wire [1:0] csr_io_pmp_7_cfg_a;
  wire  csr_io_pmp_7_cfg_x;
  wire  csr_io_pmp_7_cfg_w;
  wire  csr_io_pmp_7_cfg_r;
  wire [29:0] csr_io_pmp_7_addr;
  wire [31:0] csr_io_pmp_7_mask;
  wire  _T_1316;
  wire  _T_1317;
  wire  _T_1318;
  wire  _T_1319;
  wire  id_csr_en;
  wire  id_system_insn;
  wire  id_csr_ren;
  wire [2:0] id_csr;
  wire  _T_1330;
  wire  id_sfence;
  wire  _T_1331;
  wire  _T_1333;
  wire  _T_1334;
  wire  _T_1335;
  wire  id_csr_flush;
  wire  _T_1337;
  wire  _T_1338;
  wire  _T_1340;
  wire  _T_1341;
  wire  _T_1342;
  wire  _T_1343;
  wire  _T_1345;
  wire  _T_1346;
  wire  _T_1347;
  wire  _T_1356;
  wire  _T_1358;
  wire  _T_1359;
  wire  _T_1360;
  wire  _T_1365;
  wire  _T_1366;
  wire  _T_1367;
  wire  _T_1368;
  wire  _T_1370;
  wire  _T_1372;
  wire  _T_1373;
  wire  id_illegal_insn;
  wire  id_amo_aq;
  wire  id_amo_rl;
  wire  _T_1374;
  wire  id_fence_next;
  wire  _T_1376;
  wire  id_mem_busy;
  wire  _T_1378;
  wire  _GEN_0;
  wire  _T_1385;
  wire  _T_1388;
  wire  _T_1389;
  wire  _T_1391;
  wire  _T_1392;
  wire  _T_1393;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_bp_0_control_action;
  wire  bpu_io_bp_0_control_chain;
  wire [1:0] bpu_io_bp_0_control_tmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_h;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_x;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_r;
  wire [31:0] bpu_io_bp_0_address;
  wire [31:0] bpu_io_pc;
  wire [31:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  bpu_io_debug_if;
  wire  bpu_io_debug_ld;
  wire  bpu_io_debug_st;
  wire  _T_1403;
  wire  _T_1404;
  wire  _T_1405;
  wire  _T_1406;
  wire  _T_1407;
  wire  _T_1408;
  wire  id_xcpt;
  wire [1:0] _T_1409;
  wire [3:0] _T_1410;
  wire [3:0] _T_1411;
  wire [3:0] _T_1412;
  wire [3:0] _T_1413;
  wire [3:0] _T_1414;
  wire [31:0] id_cause;
  wire [4:0] ex_waddr;
  wire [4:0] mem_waddr;
  wire [4:0] wb_waddr;
  wire  _T_1417;
  wire  _T_1418;
  wire  _T_1420;
  wire  _T_1421;
  wire  _T_1423;
  wire  _T_1424;
  wire  id_bypass_src_0_1;
  wire  _T_1425;
  wire  id_bypass_src_0_2;
  wire  id_bypass_src_0_3;
  wire  _T_1427;
  wire  _T_1428;
  wire  id_bypass_src_1_1;
  wire  _T_1429;
  wire  id_bypass_src_1_2;
  wire  id_bypass_src_1_3;
  reg  ex_reg_rs_bypass_0;
  reg [31:0] _RAND_77;
  reg  ex_reg_rs_bypass_1;
  reg [31:0] _RAND_78;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [31:0] _RAND_79;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [31:0] _RAND_80;
  reg [29:0] ex_reg_rs_msb_0;
  reg [31:0] _RAND_81;
  reg [29:0] ex_reg_rs_msb_1;
  reg [31:0] _RAND_82;
  wire  _T_1453;
  wire [31:0] _T_1454;
  wire  _T_1456;
  wire [31:0] _T_1457;
  wire  _T_1459;
  wire [31:0] _T_1460;
  wire [31:0] _T_1461;
  wire [31:0] ex_rs_0;
  wire  _T_1463;
  wire [31:0] _T_1464;
  wire  _T_1466;
  wire [31:0] _T_1467;
  wire  _T_1469;
  wire [31:0] _T_1470;
  wire [31:0] _T_1471;
  wire [31:0] ex_rs_1;
  wire  _T_1473;
  wire  _T_1475;
  wire  _T_1476;
  wire  _T_1477;
  wire  _T_1479;
  wire [10:0] _T_1480;
  wire [10:0] _T_1481;
  wire [10:0] _T_1482;
  wire  _T_1484;
  wire  _T_1486;
  wire  _T_1487;
  wire [7:0] _T_1488;
  wire [7:0] _T_1489;
  wire [7:0] _T_1490;
  wire  _T_1495;
  wire  _T_1498;
  wire  _T_1499;
  wire  _T_1500;
  wire  _T_1502;
  wire  _T_1503;
  wire  _T_1504;
  wire  _T_1505;
  wire  _T_1506;
  wire  _T_1507;
  wire [5:0] _T_1514;
  wire [5:0] _T_1515;
  wire  _T_1520;
  wire  _T_1523;
  wire [3:0] _T_1524;
  wire [3:0] _T_1527;
  wire [3:0] _T_1528;
  wire [3:0] _T_1529;
  wire [3:0] _T_1530;
  wire [3:0] _T_1531;
  wire  _T_1536;
  wire  _T_1540;
  wire  _T_1542;
  wire  _T_1543;
  wire  _T_1544;
  wire [9:0] _T_1545;
  wire [10:0] _T_1546;
  wire  _T_1547;
  wire [7:0] _T_1548;
  wire [8:0] _T_1549;
  wire [10:0] _T_1550;
  wire  _T_1551;
  wire [11:0] _T_1552;
  wire [20:0] _T_1553;
  wire [31:0] _T_1554;
  wire [31:0] ex_imm;
  wire [31:0] _T_1557;
  wire [31:0] _T_1559;
  wire  _T_1560;
  wire [31:0] _T_1561;
  wire  _T_1562;
  wire [31:0] ex_op1;
  wire [31:0] _T_1565;
  wire [3:0] _T_1570;
  wire  _T_1571;
  wire [3:0] _T_1572;
  wire  _T_1573;
  wire [31:0] _T_1574;
  wire  _T_1575;
  wire [31:0] ex_op2;
  wire [3:0] alu_io_fn;
  wire [31:0] alu_io_in2;
  wire [31:0] alu_io_in1;
  wire [31:0] alu_io_out;
  wire [31:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire [31:0] _T_1576;
  wire [31:0] _T_1577;
  wire  div_clock;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire [31:0] div_io_req_bits_in1;
  wire [31:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [31:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  _T_1578;
  wire  _T_1580;
  wire  _T_1582;
  wire  _T_1583;
  wire  _T_1584;
  wire  _T_1587;
  wire  _T_1591;
  wire  _GEN_1;
  wire [1:0] _T_1599;
  wire  _T_1601;
  wire [1:0] _GEN_2;
  wire [1:0] _GEN_3;
  wire  _GEN_4;
  wire [1:0] _T_1605;
  wire  _T_1607;
  wire  _T_1608;
  wire [1:0] _GEN_5;
  wire [1:0] _GEN_6;
  wire [3:0] _GEN_7;
  wire [1:0] _GEN_9;
  wire [1:0] _GEN_10;
  wire  _GEN_11;
  wire  _T_1611;
  wire  _T_1613;
  wire  _T_1615;
  wire [1:0] _T_1616;
  wire [2:0] _GEN_12;
  wire  _T_1617;
  wire  _T_1618;
  wire  _T_1619;
  wire [1:0] _T_1624;
  wire [1:0] _T_1625;
  wire [1:0] _T_1626;
  wire  _T_1628;
  wire  _T_1629;
  wire [1:0] _T_1630;
  wire [29:0] _T_1631;
  wire [1:0] _GEN_13;
  wire [29:0] _GEN_14;
  wire  _T_1632;
  wire  _T_1633;
  wire  _T_1634;
  wire [1:0] _T_1639;
  wire [1:0] _T_1640;
  wire [1:0] _T_1641;
  wire  _T_1643;
  wire  _T_1644;
  wire [1:0] _T_1645;
  wire [29:0] _T_1646;
  wire [1:0] _GEN_15;
  wire [29:0] _GEN_16;
  wire [15:0] _T_1647;
  wire [31:0] _T_1648;
  wire [1:0] _T_1650;
  wire [29:0] _T_1651;
  wire  _GEN_17;
  wire [1:0] _GEN_18;
  wire [29:0] _GEN_19;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire [1:0] _GEN_28;
  wire [1:0] _GEN_29;
  wire [2:0] _GEN_30;
  wire [3:0] _GEN_32;
  wire  _GEN_33;
  wire [4:0] _GEN_34;
  wire [2:0] _GEN_35;
  wire  _GEN_39;
  wire  _GEN_40;
  wire  _GEN_41;
  wire [2:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire  _GEN_50;
  wire  _GEN_51;
  wire [1:0] _GEN_52;
  wire [29:0] _GEN_53;
  wire  _GEN_54;
  wire [1:0] _GEN_55;
  wire [29:0] _GEN_56;
  wire  _T_1654;
  wire  _T_1655;
  wire [31:0] _GEN_57;
  wire [31:0] _GEN_58;
  wire [31:0] _GEN_59;
  wire  _T_1656;
  wire  ex_pc_valid;
  wire  _T_1658;
  wire  wb_dcache_miss;
  wire  _T_1660;
  wire  _T_1661;
  wire  _T_1663;
  wire  _T_1664;
  wire  replay_ex_structural;
  wire  replay_ex_load_use;
  wire  _T_1665;
  wire  _T_1666;
  wire  replay_ex;
  wire  _T_1667;
  wire  _T_1669;
  wire  ctrl_killx;
  wire  _T_1671;
  wire  _T_1685;
  wire  _T_1686;
  wire  _T_1687;
  wire  _T_1688;
  wire  _T_1691;
  wire  _T_1692;
  wire  _T_1693;
  wire  ex_slow_bypass;
  wire  ex_xcpt;
  wire  _T_1698;
  wire  mem_pc_valid;
  wire  mem_br_taken;
  wire [31:0] _T_1699;
  wire  _T_1700;
  wire  _T_1705;
  wire  _T_1706;
  wire [10:0] _T_1712;
  wire [7:0] _T_1718;
  wire [7:0] _T_1719;
  wire [7:0] _T_1720;
  wire  _T_1729;
  wire  _T_1730;
  wire  _T_1733;
  wire  _T_1734;
  wire [5:0] _T_1744;
  wire [3:0] _T_1754;
  wire [3:0] _T_1758;
  wire [9:0] _T_1775;
  wire [10:0] _T_1776;
  wire  _T_1777;
  wire [7:0] _T_1778;
  wire [8:0] _T_1779;
  wire [10:0] _T_1780;
  wire  _T_1781;
  wire [11:0] _T_1782;
  wire [20:0] _T_1783;
  wire [31:0] _T_1784;
  wire [31:0] _T_1785;
  wire [9:0] _T_1860;
  wire [10:0] _T_1861;
  wire  _T_1862;
  wire [7:0] _T_1863;
  wire [8:0] _T_1864;
  wire [20:0] _T_1868;
  wire [31:0] _T_1869;
  wire [31:0] _T_1870;
  wire [3:0] _T_1873;
  wire [31:0] _T_1874;
  wire [31:0] _T_1875;
  wire [32:0] _T_1876;
  wire [31:0] _T_1877;
  wire [31:0] mem_br_target;
  wire  _T_1878;
  wire [31:0] _T_1879;
  wire [31:0] _T_1880;
  wire [31:0] _T_1882;
  wire [31:0] _T_1883;
  wire [31:0] mem_npc;
  wire  _T_1892;
  wire  _T_1893;
  wire  _T_1895;
  wire  mem_npc_misaligned;
  wire  _T_1897;
  wire  _T_1898;
  wire  _T_1899;
  wire [31:0] _T_1901;
  wire [31:0] mem_int_wdata;
  wire  _T_1904;
  wire  mem_cfi_taken;
  wire  _T_1909;
  wire  _T_1910;
  wire  _T_1911;
  wire  _T_1912;
  wire  _T_1914;
  wire  _T_1917;
  wire  _T_1920;
  wire  _T_1923;
  wire  _T_1925;
  wire  _T_1927;
  wire  _T_1928;
  wire  _T_1931;
  wire  _T_1936;
  wire  _T_1937;
  wire  _T_1938;
  wire  _T_1939;
  wire  _T_1940;
  wire  _T_1941;
  wire  _T_1942;
  wire  _T_1948;
  wire  _T_1949;
  wire  _T_1950;
  wire  _T_1951;
  wire  _T_1952;
  wire  _T_1953;
  wire  _T_1954;
  wire  _T_1955;
  wire  _T_1956;
  wire  _T_1957;
  wire  _T_1958;
  wire  _T_1959;
  wire  _T_1961;
  wire  _T_1963;
  wire  _T_1964;
  wire  _T_1967;
  wire  _T_1994;
  wire  _T_1995;
  wire  _T_1996;
  wire  _T_1998;
  wire [2:0] _T_2000;
  wire [1:0] _T_2002;
  wire  _T_2004;
  wire [7:0] _T_2005;
  wire [15:0] _T_2006;
  wire [31:0] _T_2007;
  wire  _T_2009;
  wire [15:0] _T_2010;
  wire [31:0] _T_2011;
  wire [31:0] _T_2012;
  wire [31:0] _T_2013;
  wire [31:0] _GEN_69;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_83;
  wire [2:0] _GEN_85;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _GEN_91;
  wire [2:0] _GEN_92;
  wire  _GEN_93;
  wire  _GEN_97;
  wire  _GEN_98;
  wire  _GEN_99;
  wire  _GEN_100;
  wire  _GEN_111;
  wire  _GEN_112;
  wire [31:0] _GEN_113;
  wire [31:0] _GEN_114;
  wire [31:0] _GEN_115;
  wire [31:0] _GEN_116;
  wire [31:0] _GEN_117;
  wire  _T_2014;
  wire  _T_2015;
  wire  mem_breakpoint;
  wire  _T_2016;
  wire  _T_2017;
  wire  mem_debug_breakpoint;
  wire  _T_2021;
  wire  mem_new_xcpt;
  wire [1:0] _T_2022;
  wire [3:0] mem_new_cause;
  wire  _T_2023;
  wire  _T_2024;
  wire  mem_xcpt;
  wire [31:0] mem_cause;
  wire  dcache_kill_mem;
  wire  _T_2026;
  wire  fpu_kill_mem;
  wire  _T_2027;
  wire  replay_mem;
  wire  _T_2028;
  wire  _T_2029;
  wire  _T_2031;
  wire  killm_common;
  wire  _T_2032;
  reg  _T_2034;
  reg [31:0] _RAND_83;
  wire  _T_2035;
  wire  _T_2036;
  wire  ctrl_killm;
  wire  _T_2038;
  wire  _T_2040;
  wire  _T_2041;
  wire  _T_2044;
  wire  _T_2047;
  wire  _T_2050;
  wire  _T_2051;
  wire [31:0] _T_2052;
  wire  _GEN_119;
  wire  _GEN_122;
  wire  _GEN_133;
  wire [2:0] _GEN_135;
  wire  _GEN_139;
  wire  _GEN_140;
  wire  _GEN_141;
  wire [2:0] _GEN_142;
  wire  _GEN_143;
  wire  _GEN_147;
  wire  _GEN_148;
  wire [31:0] _GEN_149;
  wire [31:0] _GEN_151;
  wire [31:0] _GEN_152;
  wire [31:0] _GEN_153;
  wire  _T_2056;
  wire  _T_2057;
  wire  _T_2060;
  wire  _T_2063;
  wire  _T_2066;
  wire  _T_2069;
  wire  _T_2072;
  wire  _T_2074;
  wire  _T_2075;
  wire  _T_2076;
  wire  _T_2077;
  wire  _T_2078;
  wire  wb_xcpt;
  wire [2:0] _T_2079;
  wire [3:0] _T_2080;
  wire [3:0] _T_2081;
  wire [3:0] _T_2082;
  wire [3:0] _T_2083;
  wire [31:0] wb_cause;
  wire  wb_wxd;
  wire  _T_2084;
  wire  wb_set_sboard;
  wire  replay_wb_common;
  wire  _T_2087;
  wire  replay_wb_rocc;
  wire  replay_wb;
  wire [2:0] _T_2091;
  wire [2:0] _T_2092;
  wire [31:0] _GEN_181;
  wire [32:0] _T_2093;
  wire [31:0] wb_npc;
  wire  _T_2094;
  wire  _T_2095;
  wire  _T_2096;
  wire  _T_2097;
  wire  dmem_resp_xpu;
  wire [4:0] dmem_resp_waddr;
  wire  dmem_resp_valid;
  wire  dmem_resp_replay;
  wire  _T_2102;
  wire [31:0] ll_wdata;
  wire  _T_2105;
  wire  _T_2107;
  wire  _GEN_154;
  wire [4:0] _GEN_155;
  wire  _GEN_156;
  wire  _T_2111;
  wire  _T_2112;
  wire  _T_2114;
  wire  wb_valid;
  wire  wb_wen;
  wire  rf_wen;
  wire [4:0] rf_waddr;
  wire  _T_2115;
  wire  _T_2117;
  wire [31:0] _T_2118;
  wire [31:0] _T_2119;
  wire [31:0] rf_wdata;
  wire  _T_2121;
  wire [4:0] _T_2123;
  wire  _T_2125;
  wire [31:0] _GEN_157;
  wire  _T_2126;
  wire [31:0] _GEN_158;
  wire [31:0] _GEN_163;
  wire [31:0] _GEN_164;
  wire  _GEN_167;
  wire [31:0] _GEN_169;
  wire [31:0] _GEN_170;
  wire [11:0] _T_2127;
  wire [11:0] _T_2128;
  wire [2:0] _T_2130;
  wire  _T_2133;
  wire  _T_2136;
  wire  _T_2138;
  wire  _T_2139;
  reg [31:0] _T_2142;
  reg [31:0] _RAND_84;
  wire [30:0] _T_2143;
  wire [31:0] _GEN_182;
  wire [31:0] _T_2144;
  wire [31:0] _T_2147;
  wire [31:0] _T_2149;
  wire [31:0] _T_2150;
  wire [31:0] _T_2151;
  wire [31:0] _GEN_171;
  wire [31:0] _T_2153;
  wire  _T_2154;
  wire  _T_2155;
  wire  _T_2156;
  wire  _T_2158;
  wire  _T_2159;
  wire  _T_2160;
  wire [31:0] _T_2161;
  wire  _T_2162;
  wire  _T_2163;
  wire  _T_2164;
  wire  _T_2166;
  wire  _T_2167;
  wire  _T_2168;
  wire [31:0] _T_2169;
  wire  _T_2170;
  wire  _T_2171;
  wire  _T_2172;
  wire  _T_2174;
  wire  _T_2175;
  wire  _T_2176;
  wire  _T_2177;
  wire  id_sboard_hazard;
  wire  _T_2178;
  wire [31:0] _T_2180;
  wire [31:0] _T_2182;
  wire [31:0] _T_2183;
  wire  _T_2184;
  wire [31:0] _GEN_172;
  wire  _T_2186;
  wire  _T_2187;
  wire  _T_2188;
  wire  _T_2189;
  wire  _T_2190;
  wire  ex_cannot_bypass;
  wire  _T_2191;
  wire  _T_2192;
  wire  _T_2193;
  wire  _T_2194;
  wire  _T_2195;
  wire  _T_2196;
  wire  _T_2197;
  wire  _T_2198;
  wire  data_hazard_ex;
  wire  _T_2200;
  wire  _T_2202;
  wire  _T_2203;
  wire  _T_2204;
  wire  _T_2206;
  wire  _T_2207;
  wire  _T_2208;
  wire  _T_2209;
  wire  fp_data_hazard_ex;
  wire  _T_2210;
  wire  _T_2211;
  wire  id_ex_hazard;
  wire  _T_2214;
  wire  _T_2215;
  wire  _T_2216;
  wire  _T_2217;
  wire  _T_2218;
  wire  mem_cannot_bypass;
  wire  _T_2219;
  wire  _T_2220;
  wire  _T_2221;
  wire  _T_2222;
  wire  _T_2223;
  wire  _T_2224;
  wire  _T_2225;
  wire  _T_2226;
  wire  data_hazard_mem;
  wire  _T_2228;
  wire  _T_2230;
  wire  _T_2231;
  wire  _T_2232;
  wire  _T_2234;
  wire  _T_2235;
  wire  _T_2236;
  wire  _T_2237;
  wire  fp_data_hazard_mem;
  wire  _T_2238;
  wire  _T_2239;
  wire  id_mem_hazard;
  wire  _T_2240;
  wire  _T_2241;
  wire  _T_2242;
  wire  _T_2243;
  wire  _T_2244;
  wire  _T_2245;
  wire  _T_2246;
  wire  _T_2247;
  wire  _T_2248;
  wire  _T_2249;
  wire  data_hazard_wb;
  wire  _T_2251;
  wire  _T_2253;
  wire  _T_2254;
  wire  _T_2255;
  wire  _T_2257;
  wire  _T_2258;
  wire  _T_2259;
  wire  _T_2260;
  wire  fp_data_hazard_wb;
  wire  _T_2261;
  wire  _T_2262;
  wire  id_wb_hazard;
  reg  dcache_blocked;
  reg [31:0] _RAND_85;
  wire  _T_2266;
  wire  _T_2267;
  wire  _T_2276;
  wire  _T_2277;
  wire  _T_2278;
  wire  _T_2279;
  wire  _T_2280;
  wire  _T_2281;
  wire  _T_2282;
  wire  _T_2285;
  wire  _T_2286;
  wire  _T_2291;
  wire  _T_2292;
  wire  _T_2294;
  wire  _T_2295;
  wire  _T_2296;
  wire  _T_2297;
  wire  _T_2298;
  wire  ctrl_stalld;
  wire  _T_2300;
  wire  _T_2301;
  wire  _T_2302;
  wire  _T_2303;
  wire  _T_2304;
  wire  _T_2307;
  wire  _T_2308;
  wire [31:0] _T_2309;
  wire [31:0] _T_2310;
  wire  _T_2311;
  wire  _T_2313;
  wire  _T_2314;
  wire  _T_2315;
  wire  _T_2316;
  wire  _T_2319;
  wire  _T_2320;
  wire  _T_2368;
  wire [5:0] ex_dcache_tag;
  wire [31:0] _T_2370;
  wire  _T_2371;
  wire [4:0] _T_2389;
  wire [4:0] _T_2390;
  wire [31:0] _T_2396;
  wire  _T_2399;
  wire  _T_2400;
  wire [4:0] _T_2402;
  reg [31:0] _T_2405;
  reg [31:0] _RAND_86;
  reg [31:0] _T_2407;
  reg [31:0] _RAND_87;
  reg [31:0] _T_2410;
  reg [31:0] _RAND_88;
  reg [31:0] _T_2412;
  reg [31:0] _RAND_89;
  wire  _T_2414;
  IBuf ibuf (
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_imem_ready(ibuf_io_imem_ready),
    .io_imem_valid(ibuf_io_imem_valid),
    .io_imem_bits_btb_valid(ibuf_io_imem_bits_btb_valid),
    .io_imem_bits_btb_bits_taken(ibuf_io_imem_bits_btb_bits_taken),
    .io_imem_bits_btb_bits_bridx(ibuf_io_imem_bits_btb_bits_bridx),
    .io_imem_bits_pc(ibuf_io_imem_bits_pc),
    .io_imem_bits_data(ibuf_io_imem_bits_data),
    .io_imem_bits_xcpt_pf_inst(ibuf_io_imem_bits_xcpt_pf_inst),
    .io_imem_bits_xcpt_ae_inst(ibuf_io_imem_bits_xcpt_ae_inst),
    .io_imem_bits_replay(ibuf_io_imem_bits_replay),
    .io_kill(ibuf_io_kill),
    .io_pc(ibuf_io_pc),
    .io_inst_0_ready(ibuf_io_inst_0_ready),
    .io_inst_0_valid(ibuf_io_inst_0_valid),
    .io_inst_0_bits_xcpt0_pf_inst(ibuf_io_inst_0_bits_xcpt0_pf_inst),
    .io_inst_0_bits_xcpt0_ae_inst(ibuf_io_inst_0_bits_xcpt0_ae_inst),
    .io_inst_0_bits_xcpt1_pf_inst(ibuf_io_inst_0_bits_xcpt1_pf_inst),
    .io_inst_0_bits_xcpt1_ae_inst(ibuf_io_inst_0_bits_xcpt1_ae_inst),
    .io_inst_0_bits_replay(ibuf_io_inst_0_bits_replay),
    .io_inst_0_bits_rvc(ibuf_io_inst_0_bits_rvc),
    .io_inst_0_bits_inst_bits(ibuf_io_inst_0_bits_inst_bits),
    .io_inst_0_bits_inst_rd(ibuf_io_inst_0_bits_inst_rd),
    .io_inst_0_bits_inst_rs1(ibuf_io_inst_0_bits_inst_rs1),
    .io_inst_0_bits_inst_rs2(ibuf_io_inst_0_bits_inst_rs2),
    .io_inst_0_bits_inst_rs3(ibuf_io_inst_0_bits_inst_rs3),
    .io_inst_0_bits_raw(ibuf_io_inst_0_bits_raw)
  );
  CSRFile csr (
    .clock(csr_clock),
    .reset(csr_reset),
    .io_interrupts_debug(csr_io_interrupts_debug),
    .io_interrupts_mtip(csr_io_interrupts_mtip),
    .io_interrupts_msip(csr_io_interrupts_msip),
    .io_interrupts_meip(csr_io_interrupts_meip),
    .io_hartid(csr_io_hartid),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_decode_csr(csr_io_decode_csr),
    .io_decode_read_illegal(csr_io_decode_read_illegal),
    .io_decode_write_illegal(csr_io_decode_write_illegal),
    .io_decode_write_flush(csr_io_decode_write_flush),
    .io_decode_system_illegal(csr_io_decode_system_illegal),
    .io_csr_stall(csr_io_csr_stall),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_isa(csr_io_status_isa),
    .io_status_dprv(csr_io_status_dprv),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_sxl(csr_io_status_sxl),
    .io_status_uxl(csr_io_status_uxl),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_time(csr_io_time),
    .io_rocc_interrupt(csr_io_rocc_interrupt),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_action(csr_io_bp_0_control_action),
    .io_bp_0_control_chain(csr_io_bp_0_control_chain),
    .io_bp_0_control_tmatch(csr_io_bp_0_control_tmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_h(csr_io_bp_0_control_h),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_address(csr_io_bp_0_address),
    .io_pmp_0_cfg_l(csr_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(csr_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(csr_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(csr_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(csr_io_pmp_0_cfg_r),
    .io_pmp_0_addr(csr_io_pmp_0_addr),
    .io_pmp_0_mask(csr_io_pmp_0_mask),
    .io_pmp_1_cfg_l(csr_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(csr_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(csr_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(csr_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(csr_io_pmp_1_cfg_r),
    .io_pmp_1_addr(csr_io_pmp_1_addr),
    .io_pmp_1_mask(csr_io_pmp_1_mask),
    .io_pmp_2_cfg_l(csr_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(csr_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(csr_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(csr_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(csr_io_pmp_2_cfg_r),
    .io_pmp_2_addr(csr_io_pmp_2_addr),
    .io_pmp_2_mask(csr_io_pmp_2_mask),
    .io_pmp_3_cfg_l(csr_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(csr_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(csr_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(csr_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(csr_io_pmp_3_cfg_r),
    .io_pmp_3_addr(csr_io_pmp_3_addr),
    .io_pmp_3_mask(csr_io_pmp_3_mask),
    .io_pmp_4_cfg_l(csr_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(csr_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(csr_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(csr_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(csr_io_pmp_4_cfg_r),
    .io_pmp_4_addr(csr_io_pmp_4_addr),
    .io_pmp_4_mask(csr_io_pmp_4_mask),
    .io_pmp_5_cfg_l(csr_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(csr_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(csr_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(csr_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(csr_io_pmp_5_cfg_r),
    .io_pmp_5_addr(csr_io_pmp_5_addr),
    .io_pmp_5_mask(csr_io_pmp_5_mask),
    .io_pmp_6_cfg_l(csr_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(csr_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(csr_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(csr_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(csr_io_pmp_6_cfg_r),
    .io_pmp_6_addr(csr_io_pmp_6_addr),
    .io_pmp_6_mask(csr_io_pmp_6_mask),
    .io_pmp_7_cfg_l(csr_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(csr_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(csr_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(csr_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(csr_io_pmp_7_cfg_r),
    .io_pmp_7_addr(csr_io_pmp_7_addr),
    .io_pmp_7_mask(csr_io_pmp_7_mask)
  );
  BreakpointUnit bpu (
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_bp_0_control_action(bpu_io_bp_0_control_action),
    .io_bp_0_control_chain(bpu_io_bp_0_control_chain),
    .io_bp_0_control_tmatch(bpu_io_bp_0_control_tmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_h(bpu_io_bp_0_control_h),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st),
    .io_debug_if(bpu_io_debug_if),
    .io_debug_ld(bpu_io_debug_ld),
    .io_debug_st(bpu_io_debug_st)
  );
  ALU alu (
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clock(div_clock),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  assign io_imem_req_valid = take_pc;
  assign io_imem_req_bits_pc = _T_2310;
  assign io_imem_req_bits_speculative = _T_2040;
  assign io_imem_sfence_valid = _T_2315;
  assign io_imem_sfence_bits_rs1 = _T_2316;
  assign io_imem_resp_ready = ibuf_io_imem_ready;
  assign io_imem_flush_icache = _T_2314;
  assign io_dmem_req_valid = _T_2368;
  assign io_dmem_req_bits_addr = alu_io_adder_out;
  assign io_dmem_req_bits_tag = {{1'd0}, ex_dcache_tag};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_s1_kill = _T_2371;
  assign io_dmem_s1_data_data = _T_2370;
  assign io_dmem_s1_data_mask = 4'h0;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_sfence_valid = io_imem_sfence_valid;
  assign io_ptw_sfence_bits_rs1 = io_imem_sfence_bits_rs1;
  assign io_ptw_status_dprv = csr_io_status_dprv;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_mxr = csr_io_status_mxr;
  assign io_ptw_status_sum = csr_io_status_sum;
  assign io_ptw_pmp_0_cfg_l = csr_io_pmp_0_cfg_l;
  assign io_ptw_pmp_0_cfg_a = csr_io_pmp_0_cfg_a;
  assign io_ptw_pmp_0_cfg_x = csr_io_pmp_0_cfg_x;
  assign io_ptw_pmp_0_cfg_w = csr_io_pmp_0_cfg_w;
  assign io_ptw_pmp_0_cfg_r = csr_io_pmp_0_cfg_r;
  assign io_ptw_pmp_0_addr = csr_io_pmp_0_addr;
  assign io_ptw_pmp_0_mask = csr_io_pmp_0_mask;
  assign io_ptw_pmp_1_cfg_l = csr_io_pmp_1_cfg_l;
  assign io_ptw_pmp_1_cfg_a = csr_io_pmp_1_cfg_a;
  assign io_ptw_pmp_1_cfg_x = csr_io_pmp_1_cfg_x;
  assign io_ptw_pmp_1_cfg_w = csr_io_pmp_1_cfg_w;
  assign io_ptw_pmp_1_cfg_r = csr_io_pmp_1_cfg_r;
  assign io_ptw_pmp_1_addr = csr_io_pmp_1_addr;
  assign io_ptw_pmp_1_mask = csr_io_pmp_1_mask;
  assign io_ptw_pmp_2_cfg_l = csr_io_pmp_2_cfg_l;
  assign io_ptw_pmp_2_cfg_a = csr_io_pmp_2_cfg_a;
  assign io_ptw_pmp_2_cfg_x = csr_io_pmp_2_cfg_x;
  assign io_ptw_pmp_2_cfg_w = csr_io_pmp_2_cfg_w;
  assign io_ptw_pmp_2_cfg_r = csr_io_pmp_2_cfg_r;
  assign io_ptw_pmp_2_addr = csr_io_pmp_2_addr;
  assign io_ptw_pmp_2_mask = csr_io_pmp_2_mask;
  assign io_ptw_pmp_3_cfg_l = csr_io_pmp_3_cfg_l;
  assign io_ptw_pmp_3_cfg_a = csr_io_pmp_3_cfg_a;
  assign io_ptw_pmp_3_cfg_x = csr_io_pmp_3_cfg_x;
  assign io_ptw_pmp_3_cfg_w = csr_io_pmp_3_cfg_w;
  assign io_ptw_pmp_3_cfg_r = csr_io_pmp_3_cfg_r;
  assign io_ptw_pmp_3_addr = csr_io_pmp_3_addr;
  assign io_ptw_pmp_3_mask = csr_io_pmp_3_mask;
  assign io_ptw_pmp_4_cfg_l = csr_io_pmp_4_cfg_l;
  assign io_ptw_pmp_4_cfg_a = csr_io_pmp_4_cfg_a;
  assign io_ptw_pmp_4_cfg_x = csr_io_pmp_4_cfg_x;
  assign io_ptw_pmp_4_cfg_w = csr_io_pmp_4_cfg_w;
  assign io_ptw_pmp_4_cfg_r = csr_io_pmp_4_cfg_r;
  assign io_ptw_pmp_4_addr = csr_io_pmp_4_addr;
  assign io_ptw_pmp_4_mask = csr_io_pmp_4_mask;
  assign io_ptw_pmp_5_cfg_l = csr_io_pmp_5_cfg_l;
  assign io_ptw_pmp_5_cfg_a = csr_io_pmp_5_cfg_a;
  assign io_ptw_pmp_5_cfg_x = csr_io_pmp_5_cfg_x;
  assign io_ptw_pmp_5_cfg_w = csr_io_pmp_5_cfg_w;
  assign io_ptw_pmp_5_cfg_r = csr_io_pmp_5_cfg_r;
  assign io_ptw_pmp_5_addr = csr_io_pmp_5_addr;
  assign io_ptw_pmp_5_mask = csr_io_pmp_5_mask;
  assign io_ptw_pmp_6_cfg_l = csr_io_pmp_6_cfg_l;
  assign io_ptw_pmp_6_cfg_a = csr_io_pmp_6_cfg_a;
  assign io_ptw_pmp_6_cfg_x = csr_io_pmp_6_cfg_x;
  assign io_ptw_pmp_6_cfg_w = csr_io_pmp_6_cfg_w;
  assign io_ptw_pmp_6_cfg_r = csr_io_pmp_6_cfg_r;
  assign io_ptw_pmp_6_addr = csr_io_pmp_6_addr;
  assign io_ptw_pmp_6_mask = csr_io_pmp_6_mask;
  assign io_ptw_pmp_7_cfg_l = csr_io_pmp_7_cfg_l;
  assign io_ptw_pmp_7_cfg_a = csr_io_pmp_7_cfg_a;
  assign io_ptw_pmp_7_cfg_x = csr_io_pmp_7_cfg_x;
  assign io_ptw_pmp_7_cfg_w = csr_io_pmp_7_cfg_w;
  assign io_ptw_pmp_7_cfg_r = csr_io_pmp_7_cfg_r;
  assign io_ptw_pmp_7_addr = csr_io_pmp_7_addr;
  assign io_ptw_pmp_7_mask = csr_io_pmp_7_mask;
  assign take_pc = _T_2096 | _T_1912;
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_imem_valid = io_imem_resp_valid;
  assign ibuf_io_imem_bits_btb_valid = io_imem_resp_bits_btb_valid;
  assign ibuf_io_imem_bits_btb_bits_taken = io_imem_resp_bits_btb_bits_taken;
  assign ibuf_io_imem_bits_btb_bits_bridx = io_imem_resp_bits_btb_bits_bridx;
  assign ibuf_io_imem_bits_pc = io_imem_resp_bits_pc;
  assign ibuf_io_imem_bits_data = io_imem_resp_bits_data;
  assign ibuf_io_imem_bits_xcpt_pf_inst = io_imem_resp_bits_xcpt_pf_inst;
  assign ibuf_io_imem_bits_xcpt_ae_inst = io_imem_resp_bits_xcpt_ae_inst;
  assign ibuf_io_imem_bits_replay = io_imem_resp_bits_replay;
  assign ibuf_io_kill = take_pc;
  assign ibuf_io_inst_0_ready = _T_2320;
  assign _T_679 = ibuf_io_inst_0_bits_inst_bits & 32'h505f;
  assign _T_681 = _T_679 == 32'h3;
  assign _T_683 = ibuf_io_inst_0_bits_inst_bits & 32'h207f;
  assign _T_685 = _T_683 == 32'h3;
  assign _T_687 = ibuf_io_inst_0_bits_inst_bits & 32'h607f;
  assign _T_689 = _T_687 == 32'hf;
  assign _T_691 = ibuf_io_inst_0_bits_inst_bits & 32'h5f;
  assign _T_693 = _T_691 == 32'h17;
  assign _T_695 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00007f;
  assign _T_697 = _T_695 == 32'h33;
  assign _T_699 = ibuf_io_inst_0_bits_inst_bits & 32'hbe00707f;
  assign _T_701 = _T_699 == 32'h33;
  assign _T_703 = ibuf_io_inst_0_bits_inst_bits & 32'h707b;
  assign _T_705 = _T_703 == 32'h63;
  assign _T_707 = ibuf_io_inst_0_bits_inst_bits & 32'h7f;
  assign _T_709 = _T_707 == 32'h6f;
  assign _T_711 = ibuf_io_inst_0_bits_inst_bits & 32'hffefffff;
  assign _T_713 = _T_711 == 32'h73;
  assign _T_715 = ibuf_io_inst_0_bits_inst_bits & 32'hfc00305f;
  assign _T_717 = _T_715 == 32'h1013;
  assign _T_721 = _T_683 == 32'h2013;
  assign _T_723 = ibuf_io_inst_0_bits_inst_bits & 32'h1800707f;
  assign _T_725 = _T_723 == 32'h202f;
  assign _T_729 = _T_683 == 32'h2073;
  assign _T_731 = ibuf_io_inst_0_bits_inst_bits & 32'hbc00707f;
  assign _T_733 = _T_731 == 32'h5013;
  assign _T_737 = _T_699 == 32'h5033;
  assign _T_739 = ibuf_io_inst_0_bits_inst_bits & 32'he800707f;
  assign _T_741 = _T_739 == 32'h800202f;
  assign _T_743 = ibuf_io_inst_0_bits_inst_bits & 32'hf9f0707f;
  assign _T_745 = _T_743 == 32'h1000202f;
  assign _T_747 = ibuf_io_inst_0_bits_inst_bits == 32'h10500073;
  assign _T_749 = ibuf_io_inst_0_bits_inst_bits == 32'h30200073;
  assign _T_751 = ibuf_io_inst_0_bits_inst_bits == 32'h7b200073;
  assign _T_753 = ibuf_io_inst_0_bits_inst_bits & 32'h603f;
  assign _T_755 = _T_753 == 32'h23;
  assign _T_757 = ibuf_io_inst_0_bits_inst_bits & 32'h306f;
  assign _T_759 = _T_757 == 32'h1063;
  assign _T_761 = ibuf_io_inst_0_bits_inst_bits & 32'h407f;
  assign _T_763 = _T_761 == 32'h4063;
  assign _T_767 = _T_757 == 32'h3;
  assign _T_770 = _T_681 | _T_685;
  assign _T_771 = _T_770 | _T_689;
  assign _T_772 = _T_771 | _T_693;
  assign _T_773 = _T_772 | _T_697;
  assign _T_774 = _T_773 | _T_701;
  assign _T_775 = _T_774 | _T_705;
  assign _T_776 = _T_775 | _T_709;
  assign _T_777 = _T_776 | _T_713;
  assign _T_778 = _T_777 | _T_717;
  assign _T_779 = _T_778 | _T_721;
  assign _T_780 = _T_779 | _T_725;
  assign _T_781 = _T_780 | _T_729;
  assign _T_782 = _T_781 | _T_733;
  assign _T_783 = _T_782 | _T_737;
  assign _T_784 = _T_783 | _T_741;
  assign _T_785 = _T_784 | _T_745;
  assign _T_786 = _T_785 | _T_747;
  assign _T_787 = _T_786 | _T_749;
  assign _T_788 = _T_787 | _T_751;
  assign _T_789 = _T_788 | _T_755;
  assign _T_790 = _T_789 | _T_759;
  assign _T_791 = _T_790 | _T_763;
  assign _T_792 = _T_791 | _T_767;
  assign _T_796 = ibuf_io_inst_0_bits_inst_bits & 32'h54;
  assign _T_798 = _T_796 == 32'h40;
  assign _T_802 = ibuf_io_inst_0_bits_inst_bits & 32'h48;
  assign _T_804 = _T_802 == 32'h48;
  assign _T_808 = ibuf_io_inst_0_bits_inst_bits & 32'h1c;
  assign _T_810 = _T_808 == 32'h4;
  assign _T_814 = ibuf_io_inst_0_bits_inst_bits & 32'h70;
  assign _T_816 = _T_814 == 32'h20;
  assign _T_818 = ibuf_io_inst_0_bits_inst_bits & 32'h64;
  assign _T_820 = _T_818 == 32'h20;
  assign _T_822 = ibuf_io_inst_0_bits_inst_bits & 32'h34;
  assign _T_824 = _T_822 == 32'h20;
  assign _T_827 = _T_816 | _T_820;
  assign _T_828 = _T_827 | _T_824;
  assign _T_830 = ibuf_io_inst_0_bits_inst_bits & 32'h4004;
  assign _T_832 = _T_830 == 32'h0;
  assign _T_834 = ibuf_io_inst_0_bits_inst_bits & 32'h44;
  assign _T_836 = _T_834 == 32'h0;
  assign _T_838 = ibuf_io_inst_0_bits_inst_bits & 32'h18;
  assign _T_840 = _T_838 == 32'h0;
  assign _T_842 = ibuf_io_inst_0_bits_inst_bits & 32'h2050;
  assign _T_844 = _T_842 == 32'h2000;
  assign _T_847 = _T_832 | _T_836;
  assign _T_848 = _T_847 | _T_840;
  assign _T_849 = _T_848 | _T_844;
  assign _T_851 = ibuf_io_inst_0_bits_inst_bits & 32'h58;
  assign _T_853 = _T_851 == 32'h0;
  assign _T_855 = ibuf_io_inst_0_bits_inst_bits & 32'h20;
  assign _T_857 = _T_855 == 32'h0;
  assign _T_859 = ibuf_io_inst_0_bits_inst_bits & 32'hc;
  assign _T_861 = _T_859 == 32'h4;
  assign _T_863 = ibuf_io_inst_0_bits_inst_bits & 32'h4050;
  assign _T_865 = _T_863 == 32'h4050;
  assign _T_868 = _T_853 | _T_857;
  assign _T_869 = _T_868 | _T_861;
  assign _T_870 = _T_869 | _T_804;
  assign _T_871 = _T_870 | _T_865;
  assign _T_875 = _T_802 == 32'h0;
  assign _T_877 = ibuf_io_inst_0_bits_inst_bits & 32'h4008;
  assign _T_879 = _T_877 == 32'h4000;
  assign _T_882 = _T_875 | _T_840;
  assign _T_883 = _T_882 | _T_879;
  assign _T_884 = {_T_883,_T_871};
  assign _T_886 = ibuf_io_inst_0_bits_inst_bits & 32'h50;
  assign _T_888 = _T_886 == 32'h0;
  assign _T_891 = _T_832 | _T_888;
  assign _T_892 = _T_891 | _T_836;
  assign _T_893 = _T_892 | _T_840;
  assign _T_895 = ibuf_io_inst_0_bits_inst_bits & 32'h24;
  assign _T_897 = _T_895 == 32'h4;
  assign _T_900 = _T_897 | _T_804;
  assign _T_901 = {_T_900,_T_893};
  assign _T_903 = ibuf_io_inst_0_bits_inst_bits & 32'h8;
  assign _T_905 = _T_903 == 32'h8;
  assign _T_909 = _T_834 == 32'h40;
  assign _T_912 = _T_905 | _T_909;
  assign _T_916 = _T_834 == 32'h4;
  assign _T_919 = _T_916 | _T_905;
  assign _T_923 = _T_895 == 32'h0;
  assign _T_925 = ibuf_io_inst_0_bits_inst_bits & 32'h14;
  assign _T_927 = _T_925 == 32'h10;
  assign _T_930 = _T_923 | _T_810;
  assign _T_931 = _T_930 | _T_927;
  assign _T_932 = {_T_931,_T_919};
  assign _T_933 = {_T_932,_T_912};
  assign _T_941 = ibuf_io_inst_0_bits_inst_bits & 32'h3054;
  assign _T_943 = _T_941 == 32'h1010;
  assign _T_945 = ibuf_io_inst_0_bits_inst_bits & 32'h1058;
  assign _T_947 = _T_945 == 32'h1040;
  assign _T_949 = ibuf_io_inst_0_bits_inst_bits & 32'h7044;
  assign _T_951 = _T_949 == 32'h7000;
  assign _T_954 = _T_943 | _T_947;
  assign _T_955 = _T_954 | _T_951;
  assign _T_957 = ibuf_io_inst_0_bits_inst_bits & 32'h4054;
  assign _T_959 = _T_957 == 32'h40;
  assign _T_961 = ibuf_io_inst_0_bits_inst_bits & 32'h3044;
  assign _T_963 = _T_961 == 32'h3000;
  assign _T_965 = ibuf_io_inst_0_bits_inst_bits & 32'h6044;
  assign _T_967 = _T_965 == 32'h6000;
  assign _T_969 = ibuf_io_inst_0_bits_inst_bits & 32'h6018;
  assign _T_971 = _T_969 == 32'h6000;
  assign _T_973 = ibuf_io_inst_0_bits_inst_bits & 32'h40003034;
  assign _T_975 = _T_973 == 32'h40000030;
  assign _T_977 = ibuf_io_inst_0_bits_inst_bits & 32'h40001054;
  assign _T_979 = _T_977 == 32'h40001010;
  assign _T_982 = _T_959 | _T_963;
  assign _T_983 = _T_982 | _T_967;
  assign _T_984 = _T_983 | _T_971;
  assign _T_985 = _T_984 | _T_975;
  assign _T_986 = _T_985 | _T_979;
  assign _T_988 = ibuf_io_inst_0_bits_inst_bits & 32'h2054;
  assign _T_990 = _T_988 == 32'h2010;
  assign _T_992 = ibuf_io_inst_0_bits_inst_bits & 32'h40004054;
  assign _T_994 = _T_992 == 32'h4010;
  assign _T_996 = ibuf_io_inst_0_bits_inst_bits & 32'h5054;
  assign _T_998 = _T_996 == 32'h4010;
  assign _T_1000 = ibuf_io_inst_0_bits_inst_bits & 32'h4058;
  assign _T_1002 = _T_1000 == 32'h4040;
  assign _T_1005 = _T_990 | _T_994;
  assign _T_1006 = _T_1005 | _T_998;
  assign _T_1007 = _T_1006 | _T_1002;
  assign _T_1009 = ibuf_io_inst_0_bits_inst_bits & 32'h6054;
  assign _T_1011 = _T_1009 == 32'h2010;
  assign _T_1013 = ibuf_io_inst_0_bits_inst_bits & 32'h40003054;
  assign _T_1015 = _T_1013 == 32'h40001010;
  assign _T_1018 = _T_1011 | _T_1002;
  assign _T_1019 = _T_1018 | _T_975;
  assign _T_1020 = _T_1019 | _T_1015;
  assign _T_1021 = {_T_986,_T_955};
  assign _T_1022 = {_T_1020,_T_1007};
  assign _T_1023 = {_T_1022,_T_1021};
  assign _T_1025 = ibuf_io_inst_0_bits_inst_bits & 32'h605f;
  assign _T_1027 = _T_1025 == 32'h3;
  assign _T_1029 = ibuf_io_inst_0_bits_inst_bits & 32'h707f;
  assign _T_1031 = _T_1029 == 32'h100f;
  assign _T_1034 = _T_1027 | _T_681;
  assign _T_1035 = _T_1034 | _T_685;
  assign _T_1036 = _T_1035 | _T_1031;
  assign _T_1037 = _T_1036 | _T_725;
  assign _T_1038 = _T_1037 | _T_741;
  assign _T_1039 = _T_1038 | _T_745;
  assign _T_1041 = ibuf_io_inst_0_bits_inst_bits & 32'h2008;
  assign _T_1043 = _T_1041 == 32'h8;
  assign _T_1045 = ibuf_io_inst_0_bits_inst_bits & 32'h28;
  assign _T_1047 = _T_1045 == 32'h20;
  assign _T_1049 = ibuf_io_inst_0_bits_inst_bits & 32'h18000020;
  assign _T_1051 = _T_1049 == 32'h18000020;
  assign _T_1053 = ibuf_io_inst_0_bits_inst_bits & 32'h20000020;
  assign _T_1055 = _T_1053 == 32'h20000020;
  assign _T_1058 = _T_1043 | _T_1047;
  assign _T_1059 = _T_1058 | _T_1051;
  assign _T_1060 = _T_1059 | _T_1055;
  assign _T_1062 = ibuf_io_inst_0_bits_inst_bits & 32'h10001008;
  assign _T_1064 = _T_1062 == 32'h10000008;
  assign _T_1066 = ibuf_io_inst_0_bits_inst_bits & 32'h40001008;
  assign _T_1068 = _T_1066 == 32'h40000008;
  assign _T_1071 = _T_1064 | _T_1068;
  assign _T_1073 = ibuf_io_inst_0_bits_inst_bits & 32'h8000008;
  assign _T_1075 = _T_1073 == 32'h8000008;
  assign _T_1077 = ibuf_io_inst_0_bits_inst_bits & 32'h10000008;
  assign _T_1079 = _T_1077 == 32'h10000008;
  assign _T_1081 = ibuf_io_inst_0_bits_inst_bits & 32'h80000008;
  assign _T_1083 = _T_1081 == 32'h80000008;
  assign _T_1086 = _T_1043 | _T_1075;
  assign _T_1087 = _T_1086 | _T_1079;
  assign _T_1088 = _T_1087 | _T_1083;
  assign _T_1090 = ibuf_io_inst_0_bits_inst_bits & 32'h18001008;
  assign _T_1092 = _T_1090 == 32'h8;
  assign _T_1096 = {_T_1071,_T_1060};
  assign _T_1097 = {1'h0,_T_1092};
  assign _T_1098 = {_T_1097,_T_1088};
  assign _T_1099 = {_T_1098,_T_1096};
  assign _T_1101 = ibuf_io_inst_0_bits_inst_bits & 32'h1000;
  assign _T_1103 = _T_1101 == 32'h1000;
  assign _T_1107 = ibuf_io_inst_0_bits_inst_bits & 32'h2000;
  assign _T_1109 = _T_1107 == 32'h2000;
  assign _T_1113 = ibuf_io_inst_0_bits_inst_bits & 32'h4000;
  assign _T_1115 = _T_1113 == 32'h4000;
  assign _T_1118 = {_T_1115,_T_1109};
  assign _T_1119 = {_T_1118,_T_1103};
  assign _T_1125 = ibuf_io_inst_0_bits_inst_bits & 32'h2000074;
  assign _T_1127 = _T_1125 == 32'h2000030;
  assign _T_1133 = _T_1045 == 32'h0;
  assign _T_1137 = _T_886 == 32'h10;
  assign _T_1139 = ibuf_io_inst_0_bits_inst_bits & 32'h1010;
  assign _T_1141 = _T_1139 == 32'h1010;
  assign _T_1145 = _T_1041 == 32'h2008;
  assign _T_1147 = ibuf_io_inst_0_bits_inst_bits & 32'h2010;
  assign _T_1149 = _T_1147 == 32'h2010;
  assign _T_1152 = _T_1133 | _T_861;
  assign _T_1153 = _T_1152 | _T_1137;
  assign _T_1154 = _T_1153 | _T_804;
  assign _T_1155 = _T_1154 | _T_1141;
  assign _T_1156 = _T_1155 | _T_1145;
  assign _T_1157 = _T_1156 | _T_1149;
  assign _T_1159 = ibuf_io_inst_0_bits_inst_bits & 32'h1050;
  assign _T_1161 = _T_1159 == 32'h1050;
  assign _T_1167 = _T_842 == 32'h2050;
  assign _T_1171 = ibuf_io_inst_0_bits_inst_bits & 32'h3050;
  assign _T_1173 = _T_1171 == 32'h50;
  assign _T_1176 = {_T_1173,_T_1167};
  assign _T_1177 = {_T_1176,_T_1161};
  assign _T_1179 = ibuf_io_inst_0_bits_inst_bits & 32'h1048;
  assign _T_1181 = _T_1179 == 32'h1008;
  assign _T_1185 = ibuf_io_inst_0_bits_inst_bits & 32'h3048;
  assign _T_1187 = _T_1185 == 32'h8;
  assign _T_1191 = ibuf_io_inst_0_bits_inst_bits & 32'h2048;
  assign _T_1193 = _T_1191 == 32'h2008;
  assign _T_1202__T_1211_addr = _T_1210;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_1202__T_1211_data = _T_1202[_T_1202__T_1211_addr];
  `else
  assign _T_1202__T_1211_data = _T_1202__T_1211_addr >= 5'h1f ? _RAND_75[31:0] : _T_1202[_T_1202__T_1211_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_1202__T_1221_addr = _T_1220;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_1202__T_1221_data = _T_1202[_T_1202__T_1221_addr];
  `else
  assign _T_1202__T_1221_data = _T_1202__T_1221_addr >= 5'h1f ? _RAND_76[31:0] : _T_1202[_T_1202__T_1221_addr];
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_1202__T_2124_data = rf_wdata;
  assign _T_1202__T_2124_addr = _T_2123;
  assign _T_1202__T_2124_mask = _GEN_167;
  assign _T_1202__T_2124_en = _GEN_167;
  assign _T_1206 = ibuf_io_inst_0_bits_inst_rs1 == 5'h0;
  assign _T_1209 = ibuf_io_inst_0_bits_inst_rs1;
  assign _T_1210 = ~ _T_1209;
  assign _T_1212 = _T_1202__T_1211_data;
  assign _T_1219 = ibuf_io_inst_0_bits_inst_rs2;
  assign _T_1220 = ~ _T_1219;
  assign _T_1222 = _T_1202__T_1221_data;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_interrupts_debug = io_interrupts_debug;
  assign csr_io_interrupts_mtip = io_interrupts_mtip;
  assign csr_io_interrupts_msip = io_interrupts_msip;
  assign csr_io_interrupts_meip = io_interrupts_meip;
  assign csr_io_hartid = io_hartid;
  assign csr_io_rw_addr = _T_2128;
  assign csr_io_rw_cmd = _T_2130;
  assign csr_io_rw_wdata = bypass_mux_2;
  assign csr_io_decode_csr = _T_2127;
  assign csr_io_exception = wb_xcpt;
  assign csr_io_retire = wb_valid;
  assign csr_io_cause = wb_cause;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_badaddr = bypass_mux_2;
  assign csr_io_rocc_interrupt = io_rocc_interrupt;
  assign _T_1316 = _T_1177 == 3'h2;
  assign _T_1317 = _T_1177 == 3'h3;
  assign _T_1318 = _T_1177 == 3'h1;
  assign _T_1319 = _T_1316 | _T_1317;
  assign id_csr_en = _T_1319 | _T_1318;
  assign id_system_insn = _T_1177 >= 3'h4;
  assign id_csr_ren = _T_1319 & _T_1206;
  assign id_csr = id_csr_ren ? 3'h5 : _T_1177;
  assign _T_1330 = _T_1099 == 5'h14;
  assign id_sfence = _T_1039 & _T_1330;
  assign _T_1331 = id_sfence | id_system_insn;
  assign _T_1333 = id_csr_ren == 1'h0;
  assign _T_1334 = id_csr_en & _T_1333;
  assign _T_1335 = _T_1334 & csr_io_decode_write_flush;
  assign id_csr_flush = _T_1331 | _T_1335;
  assign _T_1337 = _T_792 == 1'h0;
  assign _T_1338 = csr_io_status_isa[12];
  assign _T_1340 = _T_1338 == 1'h0;
  assign _T_1341 = _T_1127 & _T_1340;
  assign _T_1342 = _T_1337 | _T_1341;
  assign _T_1343 = csr_io_status_isa[0];
  assign _T_1345 = _T_1343 == 1'h0;
  assign _T_1346 = _T_1193 & _T_1345;
  assign _T_1347 = _T_1342 | _T_1346;
  assign _T_1356 = csr_io_status_isa[2];
  assign _T_1358 = _T_1356 == 1'h0;
  assign _T_1359 = ibuf_io_inst_0_bits_rvc & _T_1358;
  assign _T_1360 = _T_1347 | _T_1359;
  assign _T_1365 = _T_1333 & csr_io_decode_write_illegal;
  assign _T_1366 = csr_io_decode_read_illegal | _T_1365;
  assign _T_1367 = id_csr_en & _T_1366;
  assign _T_1368 = _T_1360 | _T_1367;
  assign _T_1370 = ibuf_io_inst_0_bits_rvc == 1'h0;
  assign _T_1372 = _T_1331 & csr_io_decode_system_illegal;
  assign _T_1373 = _T_1370 & _T_1372;
  assign id_illegal_insn = _T_1368 | _T_1373;
  assign id_amo_aq = ibuf_io_inst_0_bits_inst_bits[26];
  assign id_amo_rl = ibuf_io_inst_0_bits_inst_bits[25];
  assign _T_1374 = _T_1193 & id_amo_rl;
  assign id_fence_next = _T_1187 | _T_1374;
  assign _T_1376 = io_dmem_ordered == 1'h0;
  assign id_mem_busy = _T_1376 | io_dmem_req_valid;
  assign _T_1378 = id_mem_busy == 1'h0;
  assign _GEN_0 = _T_1378 ? 1'h0 : id_reg_fence;
  assign _T_1385 = wb_reg_valid & wb_ctrl_rocc;
  assign _T_1388 = _T_1193 & id_amo_aq;
  assign _T_1389 = _T_1388 | _T_1181;
  assign _T_1391 = id_reg_fence & _T_1039;
  assign _T_1392 = _T_1389 | _T_1391;
  assign _T_1393 = id_mem_busy & _T_1392;
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_bp_0_control_action = csr_io_bp_0_control_action;
  assign bpu_io_bp_0_control_chain = csr_io_bp_0_control_chain;
  assign bpu_io_bp_0_control_tmatch = csr_io_bp_0_control_tmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_h = csr_io_bp_0_control_h;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_pc = ibuf_io_pc;
  assign bpu_io_ea = bypass_mux_1;
  assign _T_1403 = csr_io_interrupt | bpu_io_debug_if;
  assign _T_1404 = _T_1403 | bpu_io_xcpt_if;
  assign _T_1405 = _T_1404 | ibuf_io_inst_0_bits_xcpt0_pf_inst;
  assign _T_1406 = _T_1405 | ibuf_io_inst_0_bits_xcpt0_ae_inst;
  assign _T_1407 = _T_1406 | ibuf_io_inst_0_bits_xcpt1_pf_inst;
  assign _T_1408 = _T_1407 | ibuf_io_inst_0_bits_xcpt1_ae_inst;
  assign id_xcpt = _T_1408 | id_illegal_insn;
  assign _T_1409 = ibuf_io_inst_0_bits_xcpt1_ae_inst ? 2'h1 : 2'h2;
  assign _T_1410 = ibuf_io_inst_0_bits_xcpt1_pf_inst ? 4'hc : {{2'd0}, _T_1409};
  assign _T_1411 = ibuf_io_inst_0_bits_xcpt0_ae_inst ? 4'h1 : _T_1410;
  assign _T_1412 = ibuf_io_inst_0_bits_xcpt0_pf_inst ? 4'hc : _T_1411;
  assign _T_1413 = bpu_io_xcpt_if ? 4'h3 : _T_1412;
  assign _T_1414 = bpu_io_debug_if ? 4'he : _T_1413;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : {{28'd0}, _T_1414};
  assign ex_waddr = ex_reg_inst[11:7];
  assign mem_waddr = mem_reg_inst[11:7];
  assign wb_waddr = wb_reg_inst[11:7];
  assign _T_1417 = ex_reg_valid & ex_ctrl_wxd;
  assign _T_1418 = mem_reg_valid & mem_ctrl_wxd;
  assign _T_1420 = mem_ctrl_mem == 1'h0;
  assign _T_1421 = _T_1418 & _T_1420;
  assign _T_1423 = 5'h0 == ibuf_io_inst_0_bits_inst_rs1;
  assign _T_1424 = ex_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign id_bypass_src_0_1 = _T_1417 & _T_1424;
  assign _T_1425 = mem_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign id_bypass_src_0_2 = _T_1421 & _T_1425;
  assign id_bypass_src_0_3 = _T_1418 & _T_1425;
  assign _T_1427 = 5'h0 == ibuf_io_inst_0_bits_inst_rs2;
  assign _T_1428 = ex_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign id_bypass_src_1_1 = _T_1417 & _T_1428;
  assign _T_1429 = mem_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign id_bypass_src_1_2 = _T_1421 & _T_1429;
  assign id_bypass_src_1_3 = _T_1418 & _T_1429;
  assign _T_1453 = ex_reg_rs_lsb_0 == 2'h1;
  assign _T_1454 = _T_1453 ? bypass_mux_1 : 32'h0;
  assign _T_1456 = ex_reg_rs_lsb_0 == 2'h2;
  assign _T_1457 = _T_1456 ? bypass_mux_2 : _T_1454;
  assign _T_1459 = ex_reg_rs_lsb_0 == 2'h3;
  assign _T_1460 = _T_1459 ? io_dmem_resp_bits_data_word_bypass : _T_1457;
  assign _T_1461 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  assign ex_rs_0 = ex_reg_rs_bypass_0 ? _T_1460 : _T_1461;
  assign _T_1463 = ex_reg_rs_lsb_1 == 2'h1;
  assign _T_1464 = _T_1463 ? bypass_mux_1 : 32'h0;
  assign _T_1466 = ex_reg_rs_lsb_1 == 2'h2;
  assign _T_1467 = _T_1466 ? bypass_mux_2 : _T_1464;
  assign _T_1469 = ex_reg_rs_lsb_1 == 2'h3;
  assign _T_1470 = _T_1469 ? io_dmem_resp_bits_data_word_bypass : _T_1467;
  assign _T_1471 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  assign ex_rs_1 = ex_reg_rs_bypass_1 ? _T_1470 : _T_1471;
  assign _T_1473 = ex_ctrl_sel_imm == 3'h5;
  assign _T_1475 = ex_reg_inst[31];
  assign _T_1476 = $signed(_T_1475);
  assign _T_1477 = _T_1473 ? $signed(1'sh0) : $signed(_T_1476);
  assign _T_1479 = ex_ctrl_sel_imm == 3'h2;
  assign _T_1480 = ex_reg_inst[30:20];
  assign _T_1481 = $signed(_T_1480);
  assign _T_1482 = _T_1479 ? $signed(_T_1481) : $signed({11{_T_1477}});
  assign _T_1484 = ex_ctrl_sel_imm != 3'h2;
  assign _T_1486 = ex_ctrl_sel_imm != 3'h3;
  assign _T_1487 = _T_1484 & _T_1486;
  assign _T_1488 = ex_reg_inst[19:12];
  assign _T_1489 = $signed(_T_1488);
  assign _T_1490 = _T_1487 ? $signed({8{_T_1477}}) : $signed(_T_1489);
  assign _T_1495 = _T_1479 | _T_1473;
  assign _T_1498 = ex_ctrl_sel_imm == 3'h3;
  assign _T_1499 = ex_reg_inst[20];
  assign _T_1500 = $signed(_T_1499);
  assign _T_1502 = ex_ctrl_sel_imm == 3'h1;
  assign _T_1503 = ex_reg_inst[7];
  assign _T_1504 = $signed(_T_1503);
  assign _T_1505 = _T_1502 ? $signed(_T_1504) : $signed(_T_1477);
  assign _T_1506 = _T_1498 ? $signed(_T_1500) : $signed(_T_1505);
  assign _T_1507 = _T_1495 ? $signed(1'sh0) : $signed(_T_1506);
  assign _T_1514 = ex_reg_inst[30:25];
  assign _T_1515 = _T_1495 ? 6'h0 : _T_1514;
  assign _T_1520 = ex_ctrl_sel_imm == 3'h0;
  assign _T_1523 = _T_1520 | _T_1502;
  assign _T_1524 = ex_reg_inst[11:8];
  assign _T_1527 = ex_reg_inst[19:16];
  assign _T_1528 = ex_reg_inst[24:21];
  assign _T_1529 = _T_1473 ? _T_1527 : _T_1528;
  assign _T_1530 = _T_1523 ? _T_1524 : _T_1529;
  assign _T_1531 = _T_1479 ? 4'h0 : _T_1530;
  assign _T_1536 = ex_ctrl_sel_imm == 3'h4;
  assign _T_1540 = ex_reg_inst[15];
  assign _T_1542 = _T_1473 ? _T_1540 : 1'h0;
  assign _T_1543 = _T_1536 ? _T_1499 : _T_1542;
  assign _T_1544 = _T_1520 ? _T_1503 : _T_1543;
  assign _T_1545 = {_T_1515,_T_1531};
  assign _T_1546 = {_T_1545,_T_1544};
  assign _T_1547 = $unsigned(_T_1507);
  assign _T_1548 = $unsigned(_T_1490);
  assign _T_1549 = {_T_1548,_T_1547};
  assign _T_1550 = $unsigned(_T_1482);
  assign _T_1551 = $unsigned(_T_1477);
  assign _T_1552 = {_T_1551,_T_1550};
  assign _T_1553 = {_T_1552,_T_1549};
  assign _T_1554 = {_T_1553,_T_1546};
  assign ex_imm = $signed(_T_1554);
  assign _T_1557 = $signed(ex_rs_0);
  assign _T_1559 = $signed(ex_reg_pc);
  assign _T_1560 = 2'h2 == ex_ctrl_sel_alu1;
  assign _T_1561 = _T_1560 ? $signed(_T_1559) : $signed(32'sh0);
  assign _T_1562 = 2'h1 == ex_ctrl_sel_alu1;
  assign ex_op1 = _T_1562 ? $signed(_T_1557) : $signed(_T_1561);
  assign _T_1565 = $signed(ex_rs_1);
  assign _T_1570 = ex_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  assign _T_1571 = 2'h1 == ex_ctrl_sel_alu2;
  assign _T_1572 = _T_1571 ? $signed(_T_1570) : $signed(4'sh0);
  assign _T_1573 = 2'h3 == ex_ctrl_sel_alu2;
  assign _T_1574 = _T_1573 ? $signed(ex_imm) : $signed({{28{_T_1572[3]}},_T_1572});
  assign _T_1575 = 2'h2 == ex_ctrl_sel_alu2;
  assign ex_op2 = _T_1575 ? $signed(_T_1565) : $signed(_T_1574);
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = _T_1576;
  assign alu_io_in1 = _T_1577;
  assign _T_1576 = $unsigned(ex_op2);
  assign _T_1577 = $unsigned(ex_op1);
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_req_valid = _T_1578;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_in1 = ex_rs_0;
  assign div_io_req_bits_in2 = ex_rs_1;
  assign div_io_req_bits_tag = ex_waddr;
  assign div_io_kill = _T_2035;
  assign div_io_resp_ready = _GEN_154;
  assign _T_1578 = ex_reg_valid & ex_ctrl_div;
  assign _T_1580 = _T_2304 == 1'h0;
  assign _T_1582 = take_pc == 1'h0;
  assign _T_1583 = _T_1582 & ibuf_io_inst_0_valid;
  assign _T_1584 = _T_1583 & ibuf_io_inst_0_bits_replay;
  assign _T_1587 = _T_1580 & id_xcpt;
  assign _T_1591 = _T_1583 & csr_io_interrupt;
  assign _GEN_1 = id_fence_next ? 1'h1 : _GEN_0;
  assign _T_1599 = {ibuf_io_inst_0_bits_xcpt1_pf_inst,ibuf_io_inst_0_bits_xcpt1_ae_inst};
  assign _T_1601 = _T_1599 != 2'h0;
  assign _GEN_2 = _T_1601 ? 2'h2 : 2'h1;
  assign _GEN_3 = _T_1601 ? 2'h1 : 2'h0;
  assign _GEN_4 = _T_1601 ? 1'h1 : ibuf_io_inst_0_bits_rvc;
  assign _T_1605 = {ibuf_io_inst_0_bits_xcpt0_pf_inst,ibuf_io_inst_0_bits_xcpt0_ae_inst};
  assign _T_1607 = _T_1605 != 2'h0;
  assign _T_1608 = bpu_io_xcpt_if | _T_1607;
  assign _GEN_5 = _T_1608 ? 2'h2 : _GEN_2;
  assign _GEN_6 = _T_1608 ? 2'h0 : _GEN_3;
  assign _GEN_7 = id_xcpt ? 4'h0 : _T_1023;
  assign _GEN_9 = id_xcpt ? _GEN_5 : _T_901;
  assign _GEN_10 = id_xcpt ? _GEN_6 : _T_884;
  assign _GEN_11 = id_xcpt ? _GEN_4 : ibuf_io_inst_0_bits_rvc;
  assign _T_1611 = _T_1181 | id_csr_flush;
  assign _T_1613 = ibuf_io_inst_0_bits_inst_rs2 != 5'h0;
  assign _T_1615 = ibuf_io_inst_0_bits_inst_rs1 != 5'h0;
  assign _T_1616 = {_T_1613,_T_1615};
  assign _GEN_12 = id_sfence ? {{1'd0}, _T_1616} : _T_1119;
  assign _T_1617 = _T_1423 | id_bypass_src_0_1;
  assign _T_1618 = _T_1617 | id_bypass_src_0_2;
  assign _T_1619 = _T_1618 | id_bypass_src_0_3;
  assign _T_1624 = id_bypass_src_0_2 ? 2'h2 : 2'h3;
  assign _T_1625 = id_bypass_src_0_1 ? 2'h1 : _T_1624;
  assign _T_1626 = _T_1423 ? 2'h0 : _T_1625;
  assign _T_1628 = _T_1619 == 1'h0;
  assign _T_1629 = _T_849 & _T_1628;
  assign _T_1630 = _GEN_169[1:0];
  assign _T_1631 = _GEN_169[31:2];
  assign _GEN_13 = _T_1629 ? _T_1630 : _T_1626;
  assign _GEN_14 = _T_1629 ? _T_1631 : ex_reg_rs_msb_0;
  assign _T_1632 = _T_1427 | id_bypass_src_1_1;
  assign _T_1633 = _T_1632 | id_bypass_src_1_2;
  assign _T_1634 = _T_1633 | id_bypass_src_1_3;
  assign _T_1639 = id_bypass_src_1_2 ? 2'h2 : 2'h3;
  assign _T_1640 = id_bypass_src_1_1 ? 2'h1 : _T_1639;
  assign _T_1641 = _T_1427 ? 2'h0 : _T_1640;
  assign _T_1643 = _T_1634 == 1'h0;
  assign _T_1644 = _T_828 & _T_1643;
  assign _T_1645 = _GEN_170[1:0];
  assign _T_1646 = _GEN_170[31:2];
  assign _GEN_15 = _T_1644 ? _T_1645 : _T_1641;
  assign _GEN_16 = _T_1644 ? _T_1646 : ex_reg_rs_msb_1;
  assign _T_1647 = ibuf_io_inst_0_bits_raw[15:0];
  assign _T_1648 = ibuf_io_inst_0_bits_rvc ? {{16'd0}, _T_1647} : ibuf_io_inst_0_bits_raw;
  assign _T_1650 = _T_1648[1:0];
  assign _T_1651 = _T_1648[31:2];
  assign _GEN_17 = id_illegal_insn ? 1'h0 : _T_1619;
  assign _GEN_18 = id_illegal_insn ? _T_1650 : _GEN_13;
  assign _GEN_19 = id_illegal_insn ? _T_1651 : _GEN_14;
  assign _GEN_21 = _T_1580 ? 1'h0 : ex_ctrl_fp;
  assign _GEN_22 = _T_1580 ? 1'h0 : ex_ctrl_rocc;
  assign _GEN_23 = _T_1580 ? _T_798 : ex_ctrl_branch;
  assign _GEN_24 = _T_1580 ? _T_804 : ex_ctrl_jal;
  assign _GEN_25 = _T_1580 ? _T_810 : ex_ctrl_jalr;
  assign _GEN_26 = _T_1580 ? _T_828 : ex_ctrl_rxs2;
  assign _GEN_28 = _T_1580 ? _GEN_10 : ex_ctrl_sel_alu2;
  assign _GEN_29 = _T_1580 ? _GEN_9 : ex_ctrl_sel_alu1;
  assign _GEN_30 = _T_1580 ? _T_933 : ex_ctrl_sel_imm;
  assign _GEN_32 = _T_1580 ? _GEN_7 : ex_ctrl_alu_fn;
  assign _GEN_33 = _T_1580 ? _T_1039 : ex_ctrl_mem;
  assign _GEN_34 = _T_1580 ? _T_1099 : ex_ctrl_mem_cmd;
  assign _GEN_35 = _T_1580 ? _GEN_12 : ex_ctrl_mem_type;
  assign _GEN_39 = _T_1580 ? 1'h0 : ex_ctrl_wfd;
  assign _GEN_40 = _T_1580 ? _T_1127 : ex_ctrl_div;
  assign _GEN_41 = _T_1580 ? _T_1157 : ex_ctrl_wxd;
  assign _GEN_42 = _T_1580 ? id_csr : ex_ctrl_csr;
  assign _GEN_43 = _T_1580 ? _T_1181 : ex_ctrl_fence_i;
  assign _GEN_47 = _T_1580 ? _GEN_11 : ex_reg_rvc;
  assign _GEN_48 = _T_1580 ? _GEN_1 : _GEN_0;
  assign _GEN_49 = _T_1580 ? _T_1611 : ex_reg_flush_pipe;
  assign _GEN_50 = _T_1580 ? _T_2241 : ex_reg_load_use;
  assign _GEN_51 = _T_1580 ? _GEN_17 : ex_reg_rs_bypass_0;
  assign _GEN_52 = _T_1580 ? _GEN_18 : ex_reg_rs_lsb_0;
  assign _GEN_53 = _T_1580 ? _GEN_19 : ex_reg_rs_msb_0;
  assign _GEN_54 = _T_1580 ? _T_1634 : ex_reg_rs_bypass_1;
  assign _GEN_55 = _T_1580 ? _GEN_15 : ex_reg_rs_lsb_1;
  assign _GEN_56 = _T_1580 ? _GEN_16 : ex_reg_rs_msb_1;
  assign _T_1654 = _T_1580 | csr_io_interrupt;
  assign _T_1655 = _T_1654 | ibuf_io_inst_0_bits_replay;
  assign _GEN_57 = _T_1655 ? id_cause : ex_cause;
  assign _GEN_58 = _T_1655 ? ibuf_io_inst_0_bits_inst_bits : ex_reg_inst;
  assign _GEN_59 = _T_1655 ? ibuf_io_pc : ex_reg_pc;
  assign _T_1656 = ex_reg_valid | ex_reg_replay;
  assign ex_pc_valid = _T_1656 | ex_reg_xcpt_interrupt;
  assign _T_1658 = io_dmem_resp_valid == 1'h0;
  assign wb_dcache_miss = wb_ctrl_mem & _T_1658;
  assign _T_1660 = io_dmem_req_ready == 1'h0;
  assign _T_1661 = ex_ctrl_mem & _T_1660;
  assign _T_1663 = div_io_req_ready == 1'h0;
  assign _T_1664 = ex_ctrl_div & _T_1663;
  assign replay_ex_structural = _T_1661 | _T_1664;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign _T_1665 = replay_ex_structural | replay_ex_load_use;
  assign _T_1666 = ex_reg_valid & _T_1665;
  assign replay_ex = ex_reg_replay | _T_1666;
  assign _T_1667 = take_pc | replay_ex;
  assign _T_1669 = ex_reg_valid == 1'h0;
  assign ctrl_killx = _T_1667 | _T_1669;
  assign _T_1671 = ex_ctrl_mem_cmd == 5'h7;
  assign _T_1685 = 3'h0 == ex_ctrl_mem_type;
  assign _T_1686 = 3'h4 == ex_ctrl_mem_type;
  assign _T_1687 = 3'h1 == ex_ctrl_mem_type;
  assign _T_1688 = 3'h5 == ex_ctrl_mem_type;
  assign _T_1691 = _T_1685 | _T_1686;
  assign _T_1692 = _T_1691 | _T_1687;
  assign _T_1693 = _T_1692 | _T_1688;
  assign ex_slow_bypass = _T_1671 | _T_1693;
  assign ex_xcpt = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign _T_1698 = mem_reg_valid | mem_reg_replay;
  assign mem_pc_valid = _T_1698 | mem_reg_xcpt_interrupt;
  assign mem_br_taken = bypass_mux_1[0];
  assign _T_1699 = $signed(mem_reg_pc);
  assign _T_1700 = mem_ctrl_branch & mem_br_taken;
  assign _T_1705 = mem_reg_inst[31];
  assign _T_1706 = $signed(_T_1705);
  assign _T_1712 = {11{_T_1706}};
  assign _T_1718 = mem_reg_inst[19:12];
  assign _T_1719 = $signed(_T_1718);
  assign _T_1720 = {8{_T_1706}};
  assign _T_1729 = mem_reg_inst[20];
  assign _T_1730 = $signed(_T_1729);
  assign _T_1733 = mem_reg_inst[7];
  assign _T_1734 = $signed(_T_1733);
  assign _T_1744 = mem_reg_inst[30:25];
  assign _T_1754 = mem_reg_inst[11:8];
  assign _T_1758 = mem_reg_inst[24:21];
  assign _T_1775 = {_T_1744,_T_1754};
  assign _T_1776 = {_T_1775,1'h0};
  assign _T_1777 = $unsigned(_T_1734);
  assign _T_1778 = $unsigned(_T_1720);
  assign _T_1779 = {_T_1778,_T_1777};
  assign _T_1780 = $unsigned(_T_1712);
  assign _T_1781 = $unsigned(_T_1706);
  assign _T_1782 = {_T_1781,_T_1780};
  assign _T_1783 = {_T_1782,_T_1779};
  assign _T_1784 = {_T_1783,_T_1776};
  assign _T_1785 = $signed(_T_1784);
  assign _T_1860 = {_T_1744,_T_1758};
  assign _T_1861 = {_T_1860,1'h0};
  assign _T_1862 = $unsigned(_T_1730);
  assign _T_1863 = $unsigned(_T_1719);
  assign _T_1864 = {_T_1863,_T_1862};
  assign _T_1868 = {_T_1782,_T_1864};
  assign _T_1869 = {_T_1868,_T_1861};
  assign _T_1870 = $signed(_T_1869);
  assign _T_1873 = mem_reg_rvc ? $signed(4'sh2) : $signed(4'sh4);
  assign _T_1874 = mem_ctrl_jal ? $signed(_T_1870) : $signed({{28{_T_1873[3]}},_T_1873});
  assign _T_1875 = _T_1700 ? $signed(_T_1785) : $signed(_T_1874);
  assign _T_1876 = $signed(_T_1699) + $signed(_T_1875);
  assign _T_1877 = _T_1876[31:0];
  assign mem_br_target = $signed(_T_1877);
  assign _T_1878 = mem_ctrl_jalr | mem_reg_sfence;
  assign _T_1879 = $signed(bypass_mux_1);
  assign _T_1880 = _T_1878 ? $signed(_T_1879) : $signed(mem_br_target);
  assign _T_1882 = $signed(_T_1880) & $signed(-32'sh2);
  assign _T_1883 = $signed(_T_1882);
  assign mem_npc = $unsigned(_T_1883);
  assign _T_1892 = mem_npc[1];
  assign _T_1893 = _T_1358 & _T_1892;
  assign _T_1895 = mem_reg_sfence == 1'h0;
  assign mem_npc_misaligned = _T_1893 & _T_1895;
  assign _T_1897 = mem_reg_xcpt == 1'h0;
  assign _T_1898 = mem_ctrl_jalr ^ mem_npc_misaligned;
  assign _T_1899 = _T_1897 & _T_1898;
  assign _T_1901 = _T_1899 ? $signed(mem_br_target) : $signed(_T_1879);
  assign mem_int_wdata = $unsigned(_T_1901);
  assign _T_1904 = _T_1700 | mem_ctrl_jalr;
  assign mem_cfi_taken = _T_1904 | mem_ctrl_jal;
  assign _T_1909 = mem_cfi_taken | mem_reg_sfence;
  assign _T_1910 = mem_ctrl_jalr & csr_io_status_debug;
  assign _T_1911 = _T_1909 | _T_1910;
  assign _T_1912 = mem_reg_valid & _T_1911;
  assign _T_1914 = ctrl_killx == 1'h0;
  assign _T_1917 = _T_1582 & replay_ex;
  assign _T_1920 = _T_1914 & ex_xcpt;
  assign _T_1923 = _T_1582 & ex_reg_xcpt_interrupt;
  assign _T_1925 = ex_ctrl_mem_cmd == 5'h0;
  assign _T_1927 = ex_ctrl_mem_cmd == 5'h6;
  assign _T_1928 = _T_1925 | _T_1927;
  assign _T_1931 = _T_1928 | _T_1671;
  assign _T_1936 = ex_ctrl_mem_cmd == 5'h4;
  assign _T_1937 = ex_ctrl_mem_cmd == 5'h9;
  assign _T_1938 = ex_ctrl_mem_cmd == 5'ha;
  assign _T_1939 = ex_ctrl_mem_cmd == 5'hb;
  assign _T_1940 = _T_1936 | _T_1937;
  assign _T_1941 = _T_1940 | _T_1938;
  assign _T_1942 = _T_1941 | _T_1939;
  assign _T_1948 = ex_ctrl_mem_cmd == 5'h8;
  assign _T_1949 = ex_ctrl_mem_cmd == 5'hc;
  assign _T_1950 = ex_ctrl_mem_cmd == 5'hd;
  assign _T_1951 = ex_ctrl_mem_cmd == 5'he;
  assign _T_1952 = ex_ctrl_mem_cmd == 5'hf;
  assign _T_1953 = _T_1948 | _T_1949;
  assign _T_1954 = _T_1953 | _T_1950;
  assign _T_1955 = _T_1954 | _T_1951;
  assign _T_1956 = _T_1955 | _T_1952;
  assign _T_1957 = _T_1942 | _T_1956;
  assign _T_1958 = _T_1931 | _T_1957;
  assign _T_1959 = ex_ctrl_mem & _T_1958;
  assign _T_1961 = ex_ctrl_mem_cmd == 5'h1;
  assign _T_1963 = ex_ctrl_mem_cmd == 5'h11;
  assign _T_1964 = _T_1961 | _T_1963;
  assign _T_1967 = _T_1964 | _T_1671;
  assign _T_1994 = _T_1967 | _T_1957;
  assign _T_1995 = ex_ctrl_mem & _T_1994;
  assign _T_1996 = ex_ctrl_mem | ex_ctrl_rocc;
  assign _T_1998 = ex_ctrl_rxs2 & _T_1996;
  assign _T_2000 = ex_ctrl_rocc ? 3'h2 : ex_ctrl_mem_type;
  assign _T_2002 = _T_2000[1:0];
  assign _T_2004 = _T_2002 == 2'h0;
  assign _T_2005 = ex_rs_1[7:0];
  assign _T_2006 = {_T_2005,_T_2005};
  assign _T_2007 = {_T_2006,_T_2006};
  assign _T_2009 = _T_2002 == 2'h1;
  assign _T_2010 = ex_rs_1[15:0];
  assign _T_2011 = {_T_2010,_T_2010};
  assign _T_2012 = _T_2009 ? _T_2011 : ex_rs_1;
  assign _T_2013 = _T_2004 ? _T_2007 : _T_2012;
  assign _GEN_69 = _T_1998 ? _T_2013 : mem_reg_rs2;
  assign _GEN_71 = ex_pc_valid ? ex_ctrl_fp : mem_ctrl_fp;
  assign _GEN_72 = ex_pc_valid ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign _GEN_73 = ex_pc_valid ? ex_ctrl_branch : mem_ctrl_branch;
  assign _GEN_74 = ex_pc_valid ? ex_ctrl_jal : mem_ctrl_jal;
  assign _GEN_75 = ex_pc_valid ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign _GEN_83 = ex_pc_valid ? ex_ctrl_mem : mem_ctrl_mem;
  assign _GEN_85 = ex_pc_valid ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign _GEN_89 = ex_pc_valid ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign _GEN_90 = ex_pc_valid ? ex_ctrl_div : mem_ctrl_div;
  assign _GEN_91 = ex_pc_valid ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign _GEN_92 = ex_pc_valid ? ex_ctrl_csr : mem_ctrl_csr;
  assign _GEN_93 = ex_pc_valid ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign _GEN_97 = ex_pc_valid ? ex_reg_rvc : mem_reg_rvc;
  assign _GEN_98 = ex_pc_valid ? _T_1959 : mem_reg_load;
  assign _GEN_99 = ex_pc_valid ? _T_1995 : mem_reg_store;
  assign _GEN_100 = ex_pc_valid ? 1'h0 : mem_reg_sfence;
  assign _GEN_111 = ex_pc_valid ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign _GEN_112 = ex_pc_valid ? ex_slow_bypass : mem_reg_slow_bypass;
  assign _GEN_113 = ex_pc_valid ? ex_cause : mem_reg_cause;
  assign _GEN_114 = ex_pc_valid ? ex_reg_inst : mem_reg_inst;
  assign _GEN_115 = ex_pc_valid ? ex_reg_pc : mem_reg_pc;
  assign _GEN_116 = ex_pc_valid ? alu_io_out : bypass_mux_1;
  assign _GEN_117 = ex_pc_valid ? _GEN_69 : mem_reg_rs2;
  assign _T_2014 = mem_reg_load & bpu_io_xcpt_ld;
  assign _T_2015 = mem_reg_store & bpu_io_xcpt_st;
  assign mem_breakpoint = _T_2014 | _T_2015;
  assign _T_2016 = mem_reg_load & bpu_io_debug_ld;
  assign _T_2017 = mem_reg_store & bpu_io_debug_st;
  assign mem_debug_breakpoint = _T_2016 | _T_2017;
  assign _T_2021 = mem_debug_breakpoint | mem_breakpoint;
  assign mem_new_xcpt = _T_2021 | mem_npc_misaligned;
  assign _T_2022 = mem_breakpoint ? 2'h3 : 2'h0;
  assign mem_new_cause = mem_debug_breakpoint ? 4'he : {{2'd0}, _T_2022};
  assign _T_2023 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign _T_2024 = mem_reg_valid & mem_new_xcpt;
  assign mem_xcpt = _T_2023 | _T_2024;
  assign mem_cause = _T_2023 ? mem_reg_cause : {{28'd0}, mem_new_cause};
  assign dcache_kill_mem = _T_1418 & io_dmem_replay_next;
  assign _T_2026 = mem_reg_valid & mem_ctrl_fp;
  assign fpu_kill_mem = _T_2026 & io_fpu_nack_mem;
  assign _T_2027 = dcache_kill_mem | mem_reg_replay;
  assign replay_mem = _T_2027 | fpu_kill_mem;
  assign _T_2028 = dcache_kill_mem | _T_2096;
  assign _T_2029 = _T_2028 | mem_reg_xcpt;
  assign _T_2031 = mem_reg_valid == 1'h0;
  assign killm_common = _T_2029 | _T_2031;
  assign _T_2032 = div_io_req_ready & div_io_req_valid;
  assign _T_2035 = killm_common & _T_2034;
  assign _T_2036 = killm_common | mem_xcpt;
  assign ctrl_killm = _T_2036 | fpu_kill_mem;
  assign _T_2038 = ctrl_killm == 1'h0;
  assign _T_2040 = _T_2096 == 1'h0;
  assign _T_2041 = replay_mem & _T_2040;
  assign _T_2044 = mem_xcpt & _T_2040;
  assign _T_2047 = _T_2038 & mem_reg_flush_pipe;
  assign _T_2050 = _T_1897 & mem_ctrl_fp;
  assign _T_2051 = _T_2050 & mem_ctrl_wxd;
  assign _T_2052 = _T_2051 ? io_fpu_toint_data : mem_int_wdata;
  assign _GEN_119 = _T_1910 ? 1'h1 : mem_ctrl_fence_i;
  assign _GEN_122 = mem_pc_valid ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign _GEN_133 = mem_pc_valid ? mem_ctrl_mem : wb_ctrl_mem;
  assign _GEN_135 = mem_pc_valid ? mem_ctrl_mem_type : wb_ctrl_mem_type;
  assign _GEN_139 = mem_pc_valid ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign _GEN_140 = mem_pc_valid ? mem_ctrl_div : wb_ctrl_div;
  assign _GEN_141 = mem_pc_valid ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign _GEN_142 = mem_pc_valid ? mem_ctrl_csr : wb_ctrl_csr;
  assign _GEN_143 = mem_pc_valid ? _GEN_119 : wb_ctrl_fence_i;
  assign _GEN_147 = mem_pc_valid ? mem_reg_rvc : wb_reg_rvc;
  assign _GEN_148 = mem_pc_valid ? mem_reg_sfence : wb_reg_sfence;
  assign _GEN_149 = mem_pc_valid ? _T_2052 : bypass_mux_2;
  assign _GEN_151 = mem_pc_valid ? mem_cause : wb_reg_cause;
  assign _GEN_152 = mem_pc_valid ? mem_reg_inst : wb_reg_inst;
  assign _GEN_153 = mem_pc_valid ? mem_reg_pc : wb_reg_pc;
  assign _T_2056 = wb_reg_valid & wb_ctrl_mem;
  assign _T_2057 = _T_2056 & io_dmem_s2_xcpt_ma_st;
  assign _T_2060 = _T_2056 & io_dmem_s2_xcpt_ma_ld;
  assign _T_2063 = _T_2056 & io_dmem_s2_xcpt_pf_st;
  assign _T_2066 = _T_2056 & io_dmem_s2_xcpt_pf_ld;
  assign _T_2069 = _T_2056 & io_dmem_s2_xcpt_ae_st;
  assign _T_2072 = _T_2056 & io_dmem_s2_xcpt_ae_ld;
  assign _T_2074 = wb_reg_xcpt | _T_2057;
  assign _T_2075 = _T_2074 | _T_2060;
  assign _T_2076 = _T_2075 | _T_2063;
  assign _T_2077 = _T_2076 | _T_2066;
  assign _T_2078 = _T_2077 | _T_2069;
  assign wb_xcpt = _T_2078 | _T_2072;
  assign _T_2079 = _T_2069 ? 3'h7 : 3'h5;
  assign _T_2080 = _T_2066 ? 4'hd : {{1'd0}, _T_2079};
  assign _T_2081 = _T_2063 ? 4'hf : _T_2080;
  assign _T_2082 = _T_2060 ? 4'h4 : _T_2081;
  assign _T_2083 = _T_2057 ? 4'h6 : _T_2082;
  assign wb_cause = wb_reg_xcpt ? wb_reg_cause : {{28'd0}, _T_2083};
  assign wb_wxd = wb_reg_valid & wb_ctrl_wxd;
  assign _T_2084 = wb_ctrl_div | wb_dcache_miss;
  assign wb_set_sboard = _T_2084 | wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  assign _T_2087 = io_rocc_cmd_ready == 1'h0;
  assign replay_wb_rocc = _T_1385 & _T_2087;
  assign replay_wb = replay_wb_common | replay_wb_rocc;
  assign _T_2091 = wb_reg_rvc ? 3'h2 : 3'h4;
  assign _T_2092 = replay_wb ? 3'h0 : _T_2091;
  assign _GEN_181 = {{29'd0}, _T_2092};
  assign _T_2093 = wb_reg_pc + _GEN_181;
  assign wb_npc = _T_2093[31:0];
  assign _T_2094 = replay_wb | wb_xcpt;
  assign _T_2095 = _T_2094 | csr_io_eret;
  assign _T_2096 = _T_2095 | wb_reg_flush_pipe;
  assign _T_2097 = io_dmem_resp_bits_tag[0];
  assign dmem_resp_xpu = _T_2097 == 1'h0;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[5:1];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  assign _T_2102 = wb_wxd == 1'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign _T_2105 = div_io_resp_ready & div_io_resp_valid;
  assign _T_2107 = dmem_resp_replay & dmem_resp_xpu;
  assign _GEN_154 = _T_2107 ? 1'h0 : _T_2102;
  assign _GEN_155 = _T_2107 ? dmem_resp_waddr : div_io_resp_bits_tag;
  assign _GEN_156 = _T_2107 ? 1'h1 : _T_2105;
  assign _T_2111 = replay_wb == 1'h0;
  assign _T_2112 = wb_reg_valid & _T_2111;
  assign _T_2114 = wb_xcpt == 1'h0;
  assign wb_valid = _T_2112 & _T_2114;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign rf_wen = wb_wen | _GEN_156;
  assign rf_waddr = _GEN_156 ? _GEN_155 : wb_waddr;
  assign _T_2115 = dmem_resp_valid & dmem_resp_xpu;
  assign _T_2117 = wb_ctrl_csr != 3'h0;
  assign _T_2118 = _T_2117 ? csr_io_rw_rdata : bypass_mux_2;
  assign _T_2119 = _GEN_156 ? ll_wdata : _T_2118;
  assign rf_wdata = _T_2115 ? io_dmem_resp_bits_data : _T_2119;
  assign _T_2121 = rf_waddr != 5'h0;
  assign _T_2123 = ~ rf_waddr;
  assign _T_2125 = rf_waddr == ibuf_io_inst_0_bits_inst_rs1;
  assign _GEN_157 = _T_2125 ? rf_wdata : _T_1212;
  assign _T_2126 = rf_waddr == ibuf_io_inst_0_bits_inst_rs2;
  assign _GEN_158 = _T_2126 ? rf_wdata : _T_1222;
  assign _GEN_163 = _T_2121 ? _GEN_157 : _T_1212;
  assign _GEN_164 = _T_2121 ? _GEN_158 : _T_1222;
  assign _GEN_167 = rf_wen ? _T_2121 : 1'h0;
  assign _GEN_169 = rf_wen ? _GEN_163 : _T_1212;
  assign _GEN_170 = rf_wen ? _GEN_164 : _T_1222;
  assign _T_2127 = ibuf_io_inst_0_bits_raw[31:20];
  assign _T_2128 = wb_reg_inst[31:20];
  assign _T_2130 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign _T_2133 = _T_849 & _T_1615;
  assign _T_2136 = _T_828 & _T_1613;
  assign _T_2138 = ibuf_io_inst_0_bits_inst_rd != 5'h0;
  assign _T_2139 = _T_1157 & _T_2138;
  assign _T_2143 = _T_2142[31:1];
  assign _GEN_182 = {{1'd0}, _T_2143};
  assign _T_2144 = _GEN_182 << 1;
  assign _T_2147 = 32'h1 << _GEN_155;
  assign _T_2149 = _GEN_156 ? _T_2147 : 32'h0;
  assign _T_2150 = ~ _T_2149;
  assign _T_2151 = _T_2144 & _T_2150;
  assign _GEN_171 = _GEN_156 ? _T_2151 : _T_2142;
  assign _T_2153 = _T_2144 >> ibuf_io_inst_0_bits_inst_rs1;
  assign _T_2154 = _T_2153[0];
  assign _T_2155 = _GEN_155 == ibuf_io_inst_0_bits_inst_rs1;
  assign _T_2156 = _GEN_156 & _T_2155;
  assign _T_2158 = _T_2156 == 1'h0;
  assign _T_2159 = _T_2154 & _T_2158;
  assign _T_2160 = _T_2133 & _T_2159;
  assign _T_2161 = _T_2144 >> ibuf_io_inst_0_bits_inst_rs2;
  assign _T_2162 = _T_2161[0];
  assign _T_2163 = _GEN_155 == ibuf_io_inst_0_bits_inst_rs2;
  assign _T_2164 = _GEN_156 & _T_2163;
  assign _T_2166 = _T_2164 == 1'h0;
  assign _T_2167 = _T_2162 & _T_2166;
  assign _T_2168 = _T_2136 & _T_2167;
  assign _T_2169 = _T_2144 >> ibuf_io_inst_0_bits_inst_rd;
  assign _T_2170 = _T_2169[0];
  assign _T_2171 = _GEN_155 == ibuf_io_inst_0_bits_inst_rd;
  assign _T_2172 = _GEN_156 & _T_2171;
  assign _T_2174 = _T_2172 == 1'h0;
  assign _T_2175 = _T_2170 & _T_2174;
  assign _T_2176 = _T_2139 & _T_2175;
  assign _T_2177 = _T_2160 | _T_2168;
  assign id_sboard_hazard = _T_2177 | _T_2176;
  assign _T_2178 = wb_set_sboard & wb_wen;
  assign _T_2180 = 32'h1 << wb_waddr;
  assign _T_2182 = _T_2178 ? _T_2180 : 32'h0;
  assign _T_2183 = _T_2151 | _T_2182;
  assign _T_2184 = _GEN_156 | _T_2178;
  assign _GEN_172 = _T_2184 ? _T_2183 : _GEN_171;
  assign _T_2186 = ex_ctrl_csr != 3'h0;
  assign _T_2187 = _T_2186 | ex_ctrl_jalr;
  assign _T_2188 = _T_2187 | ex_ctrl_mem;
  assign _T_2189 = _T_2188 | ex_ctrl_div;
  assign _T_2190 = _T_2189 | ex_ctrl_fp;
  assign ex_cannot_bypass = _T_2190 | ex_ctrl_rocc;
  assign _T_2191 = ibuf_io_inst_0_bits_inst_rs1 == ex_waddr;
  assign _T_2192 = _T_2133 & _T_2191;
  assign _T_2193 = ibuf_io_inst_0_bits_inst_rs2 == ex_waddr;
  assign _T_2194 = _T_2136 & _T_2193;
  assign _T_2195 = ibuf_io_inst_0_bits_inst_rd == ex_waddr;
  assign _T_2196 = _T_2139 & _T_2195;
  assign _T_2197 = _T_2192 | _T_2194;
  assign _T_2198 = _T_2197 | _T_2196;
  assign data_hazard_ex = ex_ctrl_wxd & _T_2198;
  assign _T_2200 = io_fpu_dec_ren1 & _T_2191;
  assign _T_2202 = io_fpu_dec_ren2 & _T_2193;
  assign _T_2203 = ibuf_io_inst_0_bits_inst_rs3 == ex_waddr;
  assign _T_2204 = io_fpu_dec_ren3 & _T_2203;
  assign _T_2206 = io_fpu_dec_wen & _T_2195;
  assign _T_2207 = _T_2200 | _T_2202;
  assign _T_2208 = _T_2207 | _T_2204;
  assign _T_2209 = _T_2208 | _T_2206;
  assign fp_data_hazard_ex = ex_ctrl_wfd & _T_2209;
  assign _T_2210 = data_hazard_ex & ex_cannot_bypass;
  assign _T_2211 = _T_2210 | fp_data_hazard_ex;
  assign id_ex_hazard = ex_reg_valid & _T_2211;
  assign _T_2214 = mem_ctrl_csr != 3'h0;
  assign _T_2215 = mem_ctrl_mem & mem_reg_slow_bypass;
  assign _T_2216 = _T_2214 | _T_2215;
  assign _T_2217 = _T_2216 | mem_ctrl_div;
  assign _T_2218 = _T_2217 | mem_ctrl_fp;
  assign mem_cannot_bypass = _T_2218 | mem_ctrl_rocc;
  assign _T_2219 = ibuf_io_inst_0_bits_inst_rs1 == mem_waddr;
  assign _T_2220 = _T_2133 & _T_2219;
  assign _T_2221 = ibuf_io_inst_0_bits_inst_rs2 == mem_waddr;
  assign _T_2222 = _T_2136 & _T_2221;
  assign _T_2223 = ibuf_io_inst_0_bits_inst_rd == mem_waddr;
  assign _T_2224 = _T_2139 & _T_2223;
  assign _T_2225 = _T_2220 | _T_2222;
  assign _T_2226 = _T_2225 | _T_2224;
  assign data_hazard_mem = mem_ctrl_wxd & _T_2226;
  assign _T_2228 = io_fpu_dec_ren1 & _T_2219;
  assign _T_2230 = io_fpu_dec_ren2 & _T_2221;
  assign _T_2231 = ibuf_io_inst_0_bits_inst_rs3 == mem_waddr;
  assign _T_2232 = io_fpu_dec_ren3 & _T_2231;
  assign _T_2234 = io_fpu_dec_wen & _T_2223;
  assign _T_2235 = _T_2228 | _T_2230;
  assign _T_2236 = _T_2235 | _T_2232;
  assign _T_2237 = _T_2236 | _T_2234;
  assign fp_data_hazard_mem = mem_ctrl_wfd & _T_2237;
  assign _T_2238 = data_hazard_mem & mem_cannot_bypass;
  assign _T_2239 = _T_2238 | fp_data_hazard_mem;
  assign id_mem_hazard = mem_reg_valid & _T_2239;
  assign _T_2240 = mem_reg_valid & data_hazard_mem;
  assign _T_2241 = _T_2240 & mem_ctrl_mem;
  assign _T_2242 = ibuf_io_inst_0_bits_inst_rs1 == wb_waddr;
  assign _T_2243 = _T_2133 & _T_2242;
  assign _T_2244 = ibuf_io_inst_0_bits_inst_rs2 == wb_waddr;
  assign _T_2245 = _T_2136 & _T_2244;
  assign _T_2246 = ibuf_io_inst_0_bits_inst_rd == wb_waddr;
  assign _T_2247 = _T_2139 & _T_2246;
  assign _T_2248 = _T_2243 | _T_2245;
  assign _T_2249 = _T_2248 | _T_2247;
  assign data_hazard_wb = wb_ctrl_wxd & _T_2249;
  assign _T_2251 = io_fpu_dec_ren1 & _T_2242;
  assign _T_2253 = io_fpu_dec_ren2 & _T_2244;
  assign _T_2254 = ibuf_io_inst_0_bits_inst_rs3 == wb_waddr;
  assign _T_2255 = io_fpu_dec_ren3 & _T_2254;
  assign _T_2257 = io_fpu_dec_wen & _T_2246;
  assign _T_2258 = _T_2251 | _T_2253;
  assign _T_2259 = _T_2258 | _T_2255;
  assign _T_2260 = _T_2259 | _T_2257;
  assign fp_data_hazard_wb = wb_ctrl_wfd & _T_2260;
  assign _T_2261 = data_hazard_wb & wb_set_sboard;
  assign _T_2262 = _T_2261 | fp_data_hazard_wb;
  assign id_wb_hazard = wb_reg_valid & _T_2262;
  assign _T_2266 = io_dmem_req_valid | dcache_blocked;
  assign _T_2267 = _T_1660 & _T_2266;
  assign _T_2276 = id_ex_hazard | id_mem_hazard;
  assign _T_2277 = _T_2276 | id_wb_hazard;
  assign _T_2278 = _T_2277 | id_sboard_hazard;
  assign _T_2279 = ex_reg_valid | mem_reg_valid;
  assign _T_2280 = _T_2279 | wb_reg_valid;
  assign _T_2281 = csr_io_singleStep & _T_2280;
  assign _T_2282 = _T_2278 | _T_2281;
  assign _T_2285 = _T_1039 & dcache_blocked;
  assign _T_2286 = _T_2282 | _T_2285;
  assign _T_2291 = div_io_resp_valid & _T_2102;
  assign _T_2292 = div_io_req_ready | _T_2291;
  assign _T_2294 = _T_2292 == 1'h0;
  assign _T_2295 = _T_2294 | div_io_req_valid;
  assign _T_2296 = _T_1127 & _T_2295;
  assign _T_2297 = _T_2286 | _T_2296;
  assign _T_2298 = _T_2297 | _T_1393;
  assign ctrl_stalld = _T_2298 | csr_io_csr_stall;
  assign _T_2300 = ibuf_io_inst_0_valid == 1'h0;
  assign _T_2301 = _T_2300 | ibuf_io_inst_0_bits_replay;
  assign _T_2302 = _T_2301 | take_pc;
  assign _T_2303 = _T_2302 | ctrl_stalld;
  assign _T_2304 = _T_2303 | csr_io_interrupt;
  assign _T_2307 = wb_xcpt | csr_io_eret;
  assign _T_2308 = replay_wb | wb_reg_flush_pipe;
  assign _T_2309 = _T_2308 ? wb_npc : mem_npc;
  assign _T_2310 = _T_2307 ? csr_io_evec : _T_2309;
  assign _T_2311 = wb_reg_valid & wb_ctrl_fence_i;
  assign _T_2313 = io_dmem_s2_nack == 1'h0;
  assign _T_2314 = _T_2311 & _T_2313;
  assign _T_2315 = wb_reg_valid & wb_reg_sfence;
  assign _T_2316 = wb_ctrl_mem_type[0];
  assign _T_2319 = ctrl_stalld == 1'h0;
  assign _T_2320 = _T_2319 | csr_io_interrupt;
  assign _T_2368 = ex_reg_valid & ex_ctrl_mem;
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  assign _T_2370 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign _T_2371 = killm_common | mem_breakpoint;
  assign _T_2389 = wb_reg_inst[19:15];
  assign _T_2390 = wb_reg_inst[24:20];
  assign _T_2396 = csr_io_time;
  assign _T_2399 = _T_2178 == 1'h0;
  assign _T_2400 = rf_wen & _T_2399;
  assign _T_2402 = _T_2400 ? rf_waddr : 5'h0;
  assign _T_2414 = reset == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ex_ctrl_fp = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  ex_ctrl_rocc = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  ex_ctrl_branch = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  ex_ctrl_jal = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  ex_ctrl_jalr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  ex_ctrl_rxs2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  ex_ctrl_sel_alu2 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  ex_ctrl_sel_alu1 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  ex_ctrl_sel_imm = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  ex_ctrl_alu_fn = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  ex_ctrl_mem = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  ex_ctrl_mem_cmd = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  ex_ctrl_mem_type = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  ex_ctrl_wfd = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  ex_ctrl_div = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  ex_ctrl_wxd = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  ex_ctrl_csr = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  ex_ctrl_fence_i = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  mem_ctrl_fp = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  mem_ctrl_rocc = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  mem_ctrl_branch = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  mem_ctrl_jal = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  mem_ctrl_jalr = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  mem_ctrl_mem = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  mem_ctrl_mem_type = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  mem_ctrl_wfd = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  mem_ctrl_div = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  mem_ctrl_wxd = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  mem_ctrl_csr = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  mem_ctrl_fence_i = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  wb_ctrl_rocc = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  wb_ctrl_mem = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  wb_ctrl_mem_type = _RAND_32[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  wb_ctrl_wfd = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  wb_ctrl_div = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  wb_ctrl_wxd = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  wb_ctrl_csr = _RAND_36[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  wb_ctrl_fence_i = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  ex_reg_xcpt_interrupt = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  ex_reg_valid = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  ex_reg_rvc = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  ex_reg_xcpt = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  ex_reg_flush_pipe = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  ex_reg_load_use = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  ex_cause = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  ex_reg_replay = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  ex_reg_pc = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  ex_reg_inst = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  mem_reg_xcpt_interrupt = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  mem_reg_valid = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  mem_reg_rvc = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  mem_reg_xcpt = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  mem_reg_replay = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  mem_reg_flush_pipe = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  mem_reg_cause = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  mem_reg_slow_bypass = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  mem_reg_load = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  mem_reg_store = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  mem_reg_sfence = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  mem_reg_pc = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  mem_reg_inst = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  bypass_mux_1 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  mem_reg_rs2 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  wb_reg_valid = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  wb_reg_rvc = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  wb_reg_xcpt = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  wb_reg_replay = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  wb_reg_flush_pipe = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  wb_reg_cause = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  wb_reg_sfence = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  wb_reg_pc = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  wb_reg_inst = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  bypass_mux_2 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  id_reg_fence = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    _T_1202[initvar] = _RAND_74[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_75 = {1{$random}};
  _RAND_76 = {1{$random}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  ex_reg_rs_bypass_0 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  ex_reg_rs_bypass_1 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  ex_reg_rs_lsb_0 = _RAND_79[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  ex_reg_rs_lsb_1 = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  ex_reg_rs_msb_0 = _RAND_81[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  ex_reg_rs_msb_1 = _RAND_82[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_2034 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_2142 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  dcache_blocked = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_2405 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_2407 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_2410 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_2412 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_1580) begin
      ex_ctrl_fp <= 1'h0;
    end
    if (_T_1580) begin
      ex_ctrl_rocc <= 1'h0;
    end
    if (_T_1580) begin
      ex_ctrl_branch <= _T_798;
    end
    if (_T_1580) begin
      ex_ctrl_jal <= _T_804;
    end
    if (_T_1580) begin
      ex_ctrl_jalr <= _T_810;
    end
    if (_T_1580) begin
      ex_ctrl_rxs2 <= _T_828;
    end
    if (_T_1580) begin
      if (id_xcpt) begin
        if (_T_1608) begin
          ex_ctrl_sel_alu2 <= 2'h0;
        end else begin
          if (_T_1601) begin
            ex_ctrl_sel_alu2 <= 2'h1;
          end else begin
            ex_ctrl_sel_alu2 <= 2'h0;
          end
        end
      end else begin
        ex_ctrl_sel_alu2 <= _T_884;
      end
    end
    if (_T_1580) begin
      if (id_xcpt) begin
        if (_T_1608) begin
          ex_ctrl_sel_alu1 <= 2'h2;
        end else begin
          if (_T_1601) begin
            ex_ctrl_sel_alu1 <= 2'h2;
          end else begin
            ex_ctrl_sel_alu1 <= 2'h1;
          end
        end
      end else begin
        ex_ctrl_sel_alu1 <= _T_901;
      end
    end
    if (_T_1580) begin
      ex_ctrl_sel_imm <= _T_933;
    end
    if (_T_1580) begin
      if (id_xcpt) begin
        ex_ctrl_alu_fn <= 4'h0;
      end else begin
        ex_ctrl_alu_fn <= _T_1023;
      end
    end
    if (_T_1580) begin
      ex_ctrl_mem <= _T_1039;
    end
    if (_T_1580) begin
      ex_ctrl_mem_cmd <= _T_1099;
    end
    if (_T_1580) begin
      if (id_sfence) begin
        ex_ctrl_mem_type <= {{1'd0}, _T_1616};
      end else begin
        ex_ctrl_mem_type <= _T_1119;
      end
    end
    if (_T_1580) begin
      ex_ctrl_wfd <= 1'h0;
    end
    if (_T_1580) begin
      ex_ctrl_div <= _T_1127;
    end
    if (_T_1580) begin
      ex_ctrl_wxd <= _T_1157;
    end
    if (_T_1580) begin
      if (id_csr_ren) begin
        ex_ctrl_csr <= 3'h5;
      end else begin
        ex_ctrl_csr <= _T_1177;
      end
    end
    if (_T_1580) begin
      ex_ctrl_fence_i <= _T_1181;
    end
    if (ex_pc_valid) begin
      mem_ctrl_fp <= ex_ctrl_fp;
    end
    if (ex_pc_valid) begin
      mem_ctrl_rocc <= ex_ctrl_rocc;
    end
    if (ex_pc_valid) begin
      mem_ctrl_branch <= ex_ctrl_branch;
    end
    if (ex_pc_valid) begin
      mem_ctrl_jal <= ex_ctrl_jal;
    end
    if (ex_pc_valid) begin
      mem_ctrl_jalr <= ex_ctrl_jalr;
    end
    if (ex_pc_valid) begin
      mem_ctrl_mem <= ex_ctrl_mem;
    end
    if (ex_pc_valid) begin
      mem_ctrl_mem_type <= ex_ctrl_mem_type;
    end
    if (ex_pc_valid) begin
      mem_ctrl_wfd <= ex_ctrl_wfd;
    end
    if (ex_pc_valid) begin
      mem_ctrl_div <= ex_ctrl_div;
    end
    if (ex_pc_valid) begin
      mem_ctrl_wxd <= ex_ctrl_wxd;
    end
    if (ex_pc_valid) begin
      mem_ctrl_csr <= ex_ctrl_csr;
    end
    if (ex_pc_valid) begin
      mem_ctrl_fence_i <= ex_ctrl_fence_i;
    end
    if (mem_pc_valid) begin
      wb_ctrl_rocc <= mem_ctrl_rocc;
    end
    if (mem_pc_valid) begin
      wb_ctrl_mem <= mem_ctrl_mem;
    end
    if (mem_pc_valid) begin
      wb_ctrl_mem_type <= mem_ctrl_mem_type;
    end
    if (mem_pc_valid) begin
      wb_ctrl_wfd <= mem_ctrl_wfd;
    end
    if (mem_pc_valid) begin
      wb_ctrl_div <= mem_ctrl_div;
    end
    if (mem_pc_valid) begin
      wb_ctrl_wxd <= mem_ctrl_wxd;
    end
    if (mem_pc_valid) begin
      wb_ctrl_csr <= mem_ctrl_csr;
    end
    if (mem_pc_valid) begin
      if (_T_1910) begin
        wb_ctrl_fence_i <= 1'h1;
      end else begin
        wb_ctrl_fence_i <= mem_ctrl_fence_i;
      end
    end
    ex_reg_xcpt_interrupt <= _T_1591;
    ex_reg_valid <= _T_1580;
    if (_T_1580) begin
      if (id_xcpt) begin
        if (_T_1601) begin
          ex_reg_rvc <= 1'h1;
        end else begin
          ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
        end
      end else begin
        ex_reg_rvc <= ibuf_io_inst_0_bits_rvc;
      end
    end
    ex_reg_xcpt <= _T_1587;
    if (_T_1580) begin
      ex_reg_flush_pipe <= _T_1611;
    end
    if (_T_1580) begin
      ex_reg_load_use <= _T_2241;
    end
    if (_T_1655) begin
      if (csr_io_interrupt) begin
        ex_cause <= csr_io_interrupt_cause;
      end else begin
        ex_cause <= {{28'd0}, _T_1414};
      end
    end
    ex_reg_replay <= _T_1584;
    if (_T_1655) begin
      ex_reg_pc <= ibuf_io_pc;
    end
    if (_T_1655) begin
      ex_reg_inst <= ibuf_io_inst_0_bits_inst_bits;
    end
    mem_reg_xcpt_interrupt <= _T_1923;
    mem_reg_valid <= _T_1914;
    if (ex_pc_valid) begin
      mem_reg_rvc <= ex_reg_rvc;
    end
    mem_reg_xcpt <= _T_1920;
    mem_reg_replay <= _T_1917;
    if (ex_pc_valid) begin
      mem_reg_flush_pipe <= ex_reg_flush_pipe;
    end
    if (ex_pc_valid) begin
      mem_reg_cause <= ex_cause;
    end
    if (ex_pc_valid) begin
      mem_reg_slow_bypass <= ex_slow_bypass;
    end
    if (ex_pc_valid) begin
      mem_reg_load <= _T_1959;
    end
    if (ex_pc_valid) begin
      mem_reg_store <= _T_1995;
    end
    if (ex_pc_valid) begin
      mem_reg_sfence <= 1'h0;
    end
    if (ex_pc_valid) begin
      mem_reg_pc <= ex_reg_pc;
    end
    if (ex_pc_valid) begin
      mem_reg_inst <= ex_reg_inst;
    end
    if (ex_pc_valid) begin
      bypass_mux_1 <= alu_io_out;
    end
    if (ex_pc_valid) begin
      if (_T_1998) begin
        if (_T_2004) begin
          mem_reg_rs2 <= _T_2007;
        end else begin
          if (_T_2009) begin
            mem_reg_rs2 <= _T_2011;
          end else begin
            if (ex_reg_rs_bypass_1) begin
              if (_T_1469) begin
                mem_reg_rs2 <= io_dmem_resp_bits_data_word_bypass;
              end else begin
                if (_T_1466) begin
                  mem_reg_rs2 <= bypass_mux_2;
                end else begin
                  if (_T_1463) begin
                    mem_reg_rs2 <= bypass_mux_1;
                  end else begin
                    mem_reg_rs2 <= 32'h0;
                  end
                end
              end
            end else begin
              mem_reg_rs2 <= _T_1471;
            end
          end
        end
      end
    end
    wb_reg_valid <= _T_2038;
    if (mem_pc_valid) begin
      wb_reg_rvc <= mem_reg_rvc;
    end
    wb_reg_xcpt <= _T_2044;
    wb_reg_replay <= _T_2041;
    wb_reg_flush_pipe <= _T_2047;
    if (mem_pc_valid) begin
      if (_T_2023) begin
        wb_reg_cause <= mem_reg_cause;
      end else begin
        wb_reg_cause <= {{28'd0}, mem_new_cause};
      end
    end
    if (mem_pc_valid) begin
      wb_reg_sfence <= mem_reg_sfence;
    end
    if (mem_pc_valid) begin
      wb_reg_pc <= mem_reg_pc;
    end
    if (mem_pc_valid) begin
      wb_reg_inst <= mem_reg_inst;
    end
    if (mem_pc_valid) begin
      if (_T_2051) begin
        bypass_mux_2 <= io_fpu_toint_data;
      end else begin
        bypass_mux_2 <= mem_int_wdata;
      end
    end
    if (reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      if (_T_1580) begin
        if (id_fence_next) begin
          id_reg_fence <= 1'h1;
        end else begin
          if (_T_1378) begin
            id_reg_fence <= 1'h0;
          end
        end
      end else begin
        if (_T_1378) begin
          id_reg_fence <= 1'h0;
        end
      end
    end
    if(_T_1202__T_2124_en & _T_1202__T_2124_mask) begin
      _T_1202[_T_1202__T_2124_addr] <= _T_1202__T_2124_data;
    end
    if (_T_1580) begin
      if (id_illegal_insn) begin
        ex_reg_rs_bypass_0 <= 1'h0;
      end else begin
        ex_reg_rs_bypass_0 <= _T_1619;
      end
    end
    if (_T_1580) begin
      ex_reg_rs_bypass_1 <= _T_1634;
    end
    if (_T_1580) begin
      if (id_illegal_insn) begin
        ex_reg_rs_lsb_0 <= _T_1650;
      end else begin
        if (_T_1629) begin
          ex_reg_rs_lsb_0 <= _T_1630;
        end else begin
          if (_T_1423) begin
            ex_reg_rs_lsb_0 <= 2'h0;
          end else begin
            if (id_bypass_src_0_1) begin
              ex_reg_rs_lsb_0 <= 2'h1;
            end else begin
              if (id_bypass_src_0_2) begin
                ex_reg_rs_lsb_0 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_0 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if (_T_1580) begin
      if (_T_1644) begin
        ex_reg_rs_lsb_1 <= _T_1645;
      end else begin
        if (_T_1427) begin
          ex_reg_rs_lsb_1 <= 2'h0;
        end else begin
          if (id_bypass_src_1_1) begin
            ex_reg_rs_lsb_1 <= 2'h1;
          end else begin
            if (id_bypass_src_1_2) begin
              ex_reg_rs_lsb_1 <= 2'h2;
            end else begin
              ex_reg_rs_lsb_1 <= 2'h3;
            end
          end
        end
      end
    end
    if (_T_1580) begin
      if (id_illegal_insn) begin
        ex_reg_rs_msb_0 <= _T_1651;
      end else begin
        if (_T_1629) begin
          ex_reg_rs_msb_0 <= _T_1631;
        end
      end
    end
    if (_T_1580) begin
      if (_T_1644) begin
        ex_reg_rs_msb_1 <= _T_1646;
      end
    end
    _T_2034 <= _T_2032;
    if (reset) begin
      _T_2142 <= 32'h0;
    end else begin
      if (_T_2184) begin
        _T_2142 <= _T_2183;
      end else begin
        if (_GEN_156) begin
          _T_2142 <= _T_2151;
        end
      end
    end
    dcache_blocked <= _T_2267;
    if (ex_reg_rs_bypass_0) begin
      if (_T_1459) begin
        _T_2405 <= io_dmem_resp_bits_data_word_bypass;
      end else begin
        if (_T_1456) begin
          _T_2405 <= bypass_mux_2;
        end else begin
          if (_T_1453) begin
            _T_2405 <= bypass_mux_1;
          end else begin
            _T_2405 <= 32'h0;
          end
        end
      end
    end else begin
      _T_2405 <= _T_1461;
    end
    _T_2407 <= _T_2405;
    if (ex_reg_rs_bypass_1) begin
      if (_T_1469) begin
        _T_2410 <= io_dmem_resp_bits_data_word_bypass;
      end else begin
        if (_T_1466) begin
          _T_2410 <= bypass_mux_2;
        end else begin
          if (_T_1463) begin
            _T_2410 <= bypass_mux_1;
          end else begin
            _T_2410 <= 32'h0;
          end
        end
      end
    end else begin
      _T_2410 <= _T_1471;
    end
    _T_2412 <= _T_2410;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2414) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n",io_hartid,_T_2396,wb_valid,wb_reg_pc,_T_2402,rf_wdata,rf_wen,_T_2389,_T_2407,_T_2390,_T_2412,wb_reg_inst,wb_reg_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module RocketTile_rocket(
  input         clock,
  input         reset,
  input         io_master_0_a_ready,
  output        io_master_0_a_valid,
  output [2:0]  io_master_0_a_bits_opcode,
  output [2:0]  io_master_0_a_bits_param,
  output [3:0]  io_master_0_a_bits_size,
  output        io_master_0_a_bits_source,
  output [31:0] io_master_0_a_bits_address,
  output [3:0]  io_master_0_a_bits_mask,
  output [31:0] io_master_0_a_bits_data,
  output        io_master_0_d_ready,
  input         io_master_0_d_valid,
  input  [2:0]  io_master_0_d_bits_opcode,
  input  [3:0]  io_master_0_d_bits_size,
  input         io_master_0_d_bits_source,
  input  [31:0] io_master_0_d_bits_data,
  input         io_master_0_d_bits_error,
  output        io_slave_0_a_ready,
  input         io_slave_0_a_valid,
  input  [2:0]  io_slave_0_a_bits_opcode,
  input  [2:0]  io_slave_0_a_bits_param,
  input  [2:0]  io_slave_0_a_bits_size,
  input  [4:0]  io_slave_0_a_bits_source,
  input  [31:0] io_slave_0_a_bits_address,
  input  [3:0]  io_slave_0_a_bits_mask,
  input  [31:0] io_slave_0_a_bits_data,
  input         io_slave_0_d_ready,
  output        io_slave_0_d_valid,
  output [2:0]  io_slave_0_d_bits_opcode,
  output [1:0]  io_slave_0_d_bits_param,
  output [2:0]  io_slave_0_d_bits_size,
  output [4:0]  io_slave_0_d_bits_source,
  output        io_slave_0_d_bits_sink,
  output [31:0] io_slave_0_d_bits_data,
  output        io_slave_0_d_bits_error,
  input         io_hartid,
  input  [31:0] io_resetVector,
  input         io_interrupts_0_0,
  input         io_interrupts_0_1,
  input         io_interrupts_0_2,
  input         io_interrupts_0_3
);
  wire  tileBus_clock;
  wire  tileBus_reset;
  wire  tileBus_io_in_1_a_ready;
  wire  tileBus_io_in_1_a_valid;
  wire [2:0] tileBus_io_in_1_a_bits_opcode;
  wire [2:0] tileBus_io_in_1_a_bits_param;
  wire [3:0] tileBus_io_in_1_a_bits_size;
  wire  tileBus_io_in_1_a_bits_source;
  wire [31:0] tileBus_io_in_1_a_bits_address;
  wire [3:0] tileBus_io_in_1_a_bits_mask;
  wire [31:0] tileBus_io_in_1_a_bits_data;
  wire  tileBus_io_in_1_d_ready;
  wire  tileBus_io_in_1_d_valid;
  wire [2:0] tileBus_io_in_1_d_bits_opcode;
  wire [3:0] tileBus_io_in_1_d_bits_size;
  wire [31:0] tileBus_io_in_1_d_bits_data;
  wire  tileBus_io_in_1_d_bits_error;
  wire  tileBus_io_in_0_a_ready;
  wire  tileBus_io_in_0_a_valid;
  wire [2:0] tileBus_io_in_0_a_bits_opcode;
  wire [2:0] tileBus_io_in_0_a_bits_param;
  wire [3:0] tileBus_io_in_0_a_bits_size;
  wire [31:0] tileBus_io_in_0_a_bits_address;
  wire [3:0] tileBus_io_in_0_a_bits_mask;
  wire [31:0] tileBus_io_in_0_a_bits_data;
  wire  tileBus_io_in_0_b_valid;
  wire [1:0] tileBus_io_in_0_b_bits_param;
  wire [31:0] tileBus_io_in_0_b_bits_address;
  wire  tileBus_io_in_0_c_ready;
  wire  tileBus_io_in_0_d_ready;
  wire  tileBus_io_in_0_d_valid;
  wire [2:0] tileBus_io_in_0_d_bits_opcode;
  wire [3:0] tileBus_io_in_0_d_bits_size;
  wire  tileBus_io_in_0_d_bits_source;
  wire [31:0] tileBus_io_in_0_d_bits_data;
  wire  tileBus_io_in_0_e_ready;
  wire  tileBus_io_out_0_a_ready;
  wire  tileBus_io_out_0_a_valid;
  wire [2:0] tileBus_io_out_0_a_bits_opcode;
  wire [2:0] tileBus_io_out_0_a_bits_param;
  wire [3:0] tileBus_io_out_0_a_bits_size;
  wire  tileBus_io_out_0_a_bits_source;
  wire [31:0] tileBus_io_out_0_a_bits_address;
  wire [3:0] tileBus_io_out_0_a_bits_mask;
  wire [31:0] tileBus_io_out_0_a_bits_data;
  wire  tileBus_io_out_0_d_ready;
  wire  tileBus_io_out_0_d_valid;
  wire [2:0] tileBus_io_out_0_d_bits_opcode;
  wire [3:0] tileBus_io_out_0_d_bits_size;
  wire  tileBus_io_out_0_d_bits_source;
  wire [31:0] tileBus_io_out_0_d_bits_data;
  wire  tileBus_io_out_0_d_bits_error;
  wire  dcache_clock;
  wire  dcache_reset;
  wire  dcache_io_cpu_req_ready;
  wire  dcache_io_cpu_req_valid;
  wire [31:0] dcache_io_cpu_req_bits_addr;
  wire [6:0] dcache_io_cpu_req_bits_tag;
  wire [4:0] dcache_io_cpu_req_bits_cmd;
  wire [2:0] dcache_io_cpu_req_bits_typ;
  wire  dcache_io_cpu_req_bits_phys;
  wire  dcache_io_cpu_s1_kill;
  wire [31:0] dcache_io_cpu_s1_data_data;
  wire [3:0] dcache_io_cpu_s1_data_mask;
  wire  dcache_io_cpu_s2_nack;
  wire  dcache_io_cpu_resp_valid;
  wire [6:0] dcache_io_cpu_resp_bits_tag;
  wire [31:0] dcache_io_cpu_resp_bits_data;
  wire  dcache_io_cpu_resp_bits_replay;
  wire  dcache_io_cpu_resp_bits_has_data;
  wire [31:0] dcache_io_cpu_resp_bits_data_word_bypass;
  wire [31:0] dcache_io_cpu_resp_bits_data_raw;
  wire  dcache_io_cpu_replay_next;
  wire  dcache_io_cpu_s2_xcpt_ma_ld;
  wire  dcache_io_cpu_s2_xcpt_ma_st;
  wire  dcache_io_cpu_s2_xcpt_pf_ld;
  wire  dcache_io_cpu_s2_xcpt_pf_st;
  wire  dcache_io_cpu_s2_xcpt_ae_ld;
  wire  dcache_io_cpu_s2_xcpt_ae_st;
  wire  dcache_io_cpu_invalidate_lr;
  wire  dcache_io_cpu_ordered;
  wire  dcache_io_ptw_req_valid;
  wire [19:0] dcache_io_ptw_req_bits_addr;
  wire  dcache_io_ptw_resp_valid;
  wire [1:0] dcache_io_ptw_status_dprv;
  wire [1:0] dcache_io_ptw_status_prv;
  wire  dcache_io_ptw_status_mxr;
  wire  dcache_io_ptw_status_sum;
  wire  dcache_io_ptw_pmp_0_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_0_cfg_a;
  wire  dcache_io_ptw_pmp_0_cfg_x;
  wire  dcache_io_ptw_pmp_0_cfg_w;
  wire  dcache_io_ptw_pmp_0_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_0_addr;
  wire [31:0] dcache_io_ptw_pmp_0_mask;
  wire  dcache_io_ptw_pmp_1_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_1_cfg_a;
  wire  dcache_io_ptw_pmp_1_cfg_x;
  wire  dcache_io_ptw_pmp_1_cfg_w;
  wire  dcache_io_ptw_pmp_1_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_1_addr;
  wire [31:0] dcache_io_ptw_pmp_1_mask;
  wire  dcache_io_ptw_pmp_2_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_2_cfg_a;
  wire  dcache_io_ptw_pmp_2_cfg_x;
  wire  dcache_io_ptw_pmp_2_cfg_w;
  wire  dcache_io_ptw_pmp_2_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_2_addr;
  wire [31:0] dcache_io_ptw_pmp_2_mask;
  wire  dcache_io_ptw_pmp_3_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_3_cfg_a;
  wire  dcache_io_ptw_pmp_3_cfg_x;
  wire  dcache_io_ptw_pmp_3_cfg_w;
  wire  dcache_io_ptw_pmp_3_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_3_addr;
  wire [31:0] dcache_io_ptw_pmp_3_mask;
  wire  dcache_io_ptw_pmp_4_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_4_cfg_a;
  wire  dcache_io_ptw_pmp_4_cfg_x;
  wire  dcache_io_ptw_pmp_4_cfg_w;
  wire  dcache_io_ptw_pmp_4_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_4_addr;
  wire [31:0] dcache_io_ptw_pmp_4_mask;
  wire  dcache_io_ptw_pmp_5_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_5_cfg_a;
  wire  dcache_io_ptw_pmp_5_cfg_x;
  wire  dcache_io_ptw_pmp_5_cfg_w;
  wire  dcache_io_ptw_pmp_5_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_5_addr;
  wire [31:0] dcache_io_ptw_pmp_5_mask;
  wire  dcache_io_ptw_pmp_6_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_6_cfg_a;
  wire  dcache_io_ptw_pmp_6_cfg_x;
  wire  dcache_io_ptw_pmp_6_cfg_w;
  wire  dcache_io_ptw_pmp_6_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_6_addr;
  wire [31:0] dcache_io_ptw_pmp_6_mask;
  wire  dcache_io_ptw_pmp_7_cfg_l;
  wire [1:0] dcache_io_ptw_pmp_7_cfg_a;
  wire  dcache_io_ptw_pmp_7_cfg_x;
  wire  dcache_io_ptw_pmp_7_cfg_w;
  wire  dcache_io_ptw_pmp_7_cfg_r;
  wire [29:0] dcache_io_ptw_pmp_7_addr;
  wire [31:0] dcache_io_ptw_pmp_7_mask;
  wire  dcache_io_mem_0_a_ready;
  wire  dcache_io_mem_0_a_valid;
  wire [2:0] dcache_io_mem_0_a_bits_opcode;
  wire [2:0] dcache_io_mem_0_a_bits_param;
  wire [3:0] dcache_io_mem_0_a_bits_size;
  wire [31:0] dcache_io_mem_0_a_bits_address;
  wire [3:0] dcache_io_mem_0_a_bits_mask;
  wire [31:0] dcache_io_mem_0_a_bits_data;
  wire  dcache_io_mem_0_b_ready;
  wire  dcache_io_mem_0_b_valid;
  wire [1:0] dcache_io_mem_0_b_bits_param;
  wire [31:0] dcache_io_mem_0_b_bits_address;
  wire  dcache_io_mem_0_c_ready;
  wire  dcache_io_mem_0_c_valid;
  wire [31:0] dcache_io_mem_0_c_bits_address;
  wire  dcache_io_mem_0_d_ready;
  wire  dcache_io_mem_0_d_valid;
  wire [2:0] dcache_io_mem_0_d_bits_opcode;
  wire [3:0] dcache_io_mem_0_d_bits_size;
  wire  dcache_io_mem_0_d_bits_source;
  wire [31:0] dcache_io_mem_0_d_bits_data;
  wire  dcache_io_mem_0_e_ready;
  wire  dcache_io_mem_0_e_valid;
  wire  frontend_clock;
  wire  frontend_reset;
  wire  frontend_io_tl_out_0_a_ready;
  wire  frontend_io_tl_out_0_a_valid;
  wire [2:0] frontend_io_tl_out_0_a_bits_opcode;
  wire [2:0] frontend_io_tl_out_0_a_bits_param;
  wire [3:0] frontend_io_tl_out_0_a_bits_size;
  wire  frontend_io_tl_out_0_a_bits_source;
  wire [31:0] frontend_io_tl_out_0_a_bits_address;
  wire [3:0] frontend_io_tl_out_0_a_bits_mask;
  wire [31:0] frontend_io_tl_out_0_a_bits_data;
  wire  frontend_io_tl_out_0_d_ready;
  wire  frontend_io_tl_out_0_d_valid;
  wire [2:0] frontend_io_tl_out_0_d_bits_opcode;
  wire [3:0] frontend_io_tl_out_0_d_bits_size;
  wire [31:0] frontend_io_tl_out_0_d_bits_data;
  wire  frontend_io_tl_out_0_d_bits_error;
  wire  frontend_io_cpu_req_valid;
  wire [31:0] frontend_io_cpu_req_bits_pc;
  wire  frontend_io_cpu_req_bits_speculative;
  wire  frontend_io_cpu_resp_ready;
  wire  frontend_io_cpu_resp_valid;
  wire  frontend_io_cpu_resp_bits_btb_valid;
  wire  frontend_io_cpu_resp_bits_btb_bits_taken;
  wire  frontend_io_cpu_resp_bits_btb_bits_bridx;
  wire [31:0] frontend_io_cpu_resp_bits_pc;
  wire [31:0] frontend_io_cpu_resp_bits_data;
  wire  frontend_io_cpu_resp_bits_xcpt_pf_inst;
  wire  frontend_io_cpu_resp_bits_xcpt_ae_inst;
  wire  frontend_io_cpu_resp_bits_replay;
  wire  frontend_io_cpu_flush_icache;
  wire [31:0] frontend_io_cpu_npc;
  wire  frontend_io_ptw_req_valid;
  wire [19:0] frontend_io_ptw_req_bits_addr;
  wire  frontend_io_ptw_resp_valid;
  wire [1:0] frontend_io_ptw_status_dprv;
  wire [1:0] frontend_io_ptw_status_prv;
  wire  frontend_io_ptw_status_mxr;
  wire  frontend_io_ptw_status_sum;
  wire  frontend_io_ptw_pmp_0_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_0_cfg_a;
  wire  frontend_io_ptw_pmp_0_cfg_x;
  wire  frontend_io_ptw_pmp_0_cfg_w;
  wire  frontend_io_ptw_pmp_0_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_0_addr;
  wire [31:0] frontend_io_ptw_pmp_0_mask;
  wire  frontend_io_ptw_pmp_1_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_1_cfg_a;
  wire  frontend_io_ptw_pmp_1_cfg_x;
  wire  frontend_io_ptw_pmp_1_cfg_w;
  wire  frontend_io_ptw_pmp_1_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_1_addr;
  wire [31:0] frontend_io_ptw_pmp_1_mask;
  wire  frontend_io_ptw_pmp_2_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_2_cfg_a;
  wire  frontend_io_ptw_pmp_2_cfg_x;
  wire  frontend_io_ptw_pmp_2_cfg_w;
  wire  frontend_io_ptw_pmp_2_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_2_addr;
  wire [31:0] frontend_io_ptw_pmp_2_mask;
  wire  frontend_io_ptw_pmp_3_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_3_cfg_a;
  wire  frontend_io_ptw_pmp_3_cfg_x;
  wire  frontend_io_ptw_pmp_3_cfg_w;
  wire  frontend_io_ptw_pmp_3_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_3_addr;
  wire [31:0] frontend_io_ptw_pmp_3_mask;
  wire  frontend_io_ptw_pmp_4_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_4_cfg_a;
  wire  frontend_io_ptw_pmp_4_cfg_x;
  wire  frontend_io_ptw_pmp_4_cfg_w;
  wire  frontend_io_ptw_pmp_4_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_4_addr;
  wire [31:0] frontend_io_ptw_pmp_4_mask;
  wire  frontend_io_ptw_pmp_5_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_5_cfg_a;
  wire  frontend_io_ptw_pmp_5_cfg_x;
  wire  frontend_io_ptw_pmp_5_cfg_w;
  wire  frontend_io_ptw_pmp_5_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_5_addr;
  wire [31:0] frontend_io_ptw_pmp_5_mask;
  wire  frontend_io_ptw_pmp_6_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_6_cfg_a;
  wire  frontend_io_ptw_pmp_6_cfg_x;
  wire  frontend_io_ptw_pmp_6_cfg_w;
  wire  frontend_io_ptw_pmp_6_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_6_addr;
  wire [31:0] frontend_io_ptw_pmp_6_mask;
  wire  frontend_io_ptw_pmp_7_cfg_l;
  wire [1:0] frontend_io_ptw_pmp_7_cfg_a;
  wire  frontend_io_ptw_pmp_7_cfg_x;
  wire  frontend_io_ptw_pmp_7_cfg_w;
  wire  frontend_io_ptw_pmp_7_cfg_r;
  wire [29:0] frontend_io_ptw_pmp_7_addr;
  wire [31:0] frontend_io_ptw_pmp_7_mask;
  wire [31:0] frontend_io_resetVector;
  wire  ScratchpadSlavePort_clock;
  wire  ScratchpadSlavePort_reset;
  wire  ScratchpadSlavePort_io_tl_in_0_a_ready;
  wire  ScratchpadSlavePort_io_tl_in_0_a_valid;
  wire [2:0] ScratchpadSlavePort_io_tl_in_0_a_bits_opcode;
  wire [2:0] ScratchpadSlavePort_io_tl_in_0_a_bits_param;
  wire [1:0] ScratchpadSlavePort_io_tl_in_0_a_bits_size;
  wire [9:0] ScratchpadSlavePort_io_tl_in_0_a_bits_source;
  wire [31:0] ScratchpadSlavePort_io_tl_in_0_a_bits_address;
  wire [3:0] ScratchpadSlavePort_io_tl_in_0_a_bits_mask;
  wire [31:0] ScratchpadSlavePort_io_tl_in_0_a_bits_data;
  wire  ScratchpadSlavePort_io_tl_in_0_d_ready;
  wire  ScratchpadSlavePort_io_tl_in_0_d_valid;
  wire [2:0] ScratchpadSlavePort_io_tl_in_0_d_bits_opcode;
  wire [1:0] ScratchpadSlavePort_io_tl_in_0_d_bits_param;
  wire [1:0] ScratchpadSlavePort_io_tl_in_0_d_bits_size;
  wire [9:0] ScratchpadSlavePort_io_tl_in_0_d_bits_source;
  wire  ScratchpadSlavePort_io_tl_in_0_d_bits_sink;
  wire [31:0] ScratchpadSlavePort_io_tl_in_0_d_bits_data;
  wire  ScratchpadSlavePort_io_tl_in_0_d_bits_error;
  wire  ScratchpadSlavePort_io_dmem_req_ready;
  wire  ScratchpadSlavePort_io_dmem_req_valid;
  wire [31:0] ScratchpadSlavePort_io_dmem_req_bits_addr;
  wire [6:0] ScratchpadSlavePort_io_dmem_req_bits_tag;
  wire [4:0] ScratchpadSlavePort_io_dmem_req_bits_cmd;
  wire [2:0] ScratchpadSlavePort_io_dmem_req_bits_typ;
  wire  ScratchpadSlavePort_io_dmem_req_bits_phys;
  wire  ScratchpadSlavePort_io_dmem_s1_kill;
  wire [31:0] ScratchpadSlavePort_io_dmem_s1_data_data;
  wire [3:0] ScratchpadSlavePort_io_dmem_s1_data_mask;
  wire  ScratchpadSlavePort_io_dmem_s2_nack;
  wire  ScratchpadSlavePort_io_dmem_resp_valid;
  wire [31:0] ScratchpadSlavePort_io_dmem_resp_bits_data_raw;
  wire  ScratchpadSlavePort_io_dmem_invalidate_lr;
  wire  TLFragmenter_clock;
  wire  TLFragmenter_reset;
  wire  TLFragmenter_io_in_0_a_ready;
  wire  TLFragmenter_io_in_0_a_valid;
  wire [2:0] TLFragmenter_io_in_0_a_bits_opcode;
  wire [2:0] TLFragmenter_io_in_0_a_bits_param;
  wire [2:0] TLFragmenter_io_in_0_a_bits_size;
  wire [4:0] TLFragmenter_io_in_0_a_bits_source;
  wire [31:0] TLFragmenter_io_in_0_a_bits_address;
  wire [3:0] TLFragmenter_io_in_0_a_bits_mask;
  wire [31:0] TLFragmenter_io_in_0_a_bits_data;
  wire  TLFragmenter_io_in_0_d_ready;
  wire  TLFragmenter_io_in_0_d_valid;
  wire [2:0] TLFragmenter_io_in_0_d_bits_opcode;
  wire [1:0] TLFragmenter_io_in_0_d_bits_param;
  wire [2:0] TLFragmenter_io_in_0_d_bits_size;
  wire [4:0] TLFragmenter_io_in_0_d_bits_source;
  wire  TLFragmenter_io_in_0_d_bits_sink;
  wire [31:0] TLFragmenter_io_in_0_d_bits_data;
  wire  TLFragmenter_io_in_0_d_bits_error;
  wire  TLFragmenter_io_out_0_a_ready;
  wire  TLFragmenter_io_out_0_a_valid;
  wire [2:0] TLFragmenter_io_out_0_a_bits_opcode;
  wire [2:0] TLFragmenter_io_out_0_a_bits_param;
  wire [1:0] TLFragmenter_io_out_0_a_bits_size;
  wire [9:0] TLFragmenter_io_out_0_a_bits_source;
  wire [31:0] TLFragmenter_io_out_0_a_bits_address;
  wire [3:0] TLFragmenter_io_out_0_a_bits_mask;
  wire [31:0] TLFragmenter_io_out_0_a_bits_data;
  wire  TLFragmenter_io_out_0_d_ready;
  wire  TLFragmenter_io_out_0_d_valid;
  wire [2:0] TLFragmenter_io_out_0_d_bits_opcode;
  wire [1:0] TLFragmenter_io_out_0_d_bits_param;
  wire [1:0] TLFragmenter_io_out_0_d_bits_size;
  wire [9:0] TLFragmenter_io_out_0_d_bits_source;
  wire  TLFragmenter_io_out_0_d_bits_sink;
  wire [31:0] TLFragmenter_io_out_0_d_bits_data;
  wire  TLFragmenter_io_out_0_d_bits_error;
  wire  dcacheArb_clock;
  wire  dcacheArb_io_requestor_0_req_ready;
  wire  dcacheArb_io_requestor_0_req_valid;
  wire [31:0] dcacheArb_io_requestor_0_req_bits_addr;
  wire [6:0] dcacheArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcacheArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcacheArb_io_requestor_0_req_bits_typ;
  wire  dcacheArb_io_requestor_0_req_bits_phys;
  wire  dcacheArb_io_requestor_0_s1_kill;
  wire [31:0] dcacheArb_io_requestor_0_s1_data_data;
  wire [3:0] dcacheArb_io_requestor_0_s1_data_mask;
  wire  dcacheArb_io_requestor_0_s2_nack;
  wire  dcacheArb_io_requestor_0_resp_valid;
  wire [31:0] dcacheArb_io_requestor_0_resp_bits_data_raw;
  wire  dcacheArb_io_requestor_0_invalidate_lr;
  wire  dcacheArb_io_requestor_1_req_ready;
  wire  dcacheArb_io_requestor_1_req_valid;
  wire [31:0] dcacheArb_io_requestor_1_req_bits_addr;
  wire [6:0] dcacheArb_io_requestor_1_req_bits_tag;
  wire [4:0] dcacheArb_io_requestor_1_req_bits_cmd;
  wire [2:0] dcacheArb_io_requestor_1_req_bits_typ;
  wire  dcacheArb_io_requestor_1_req_bits_phys;
  wire  dcacheArb_io_requestor_1_s1_kill;
  wire [31:0] dcacheArb_io_requestor_1_s1_data_data;
  wire [3:0] dcacheArb_io_requestor_1_s1_data_mask;
  wire  dcacheArb_io_requestor_1_s2_nack;
  wire  dcacheArb_io_requestor_1_resp_valid;
  wire [6:0] dcacheArb_io_requestor_1_resp_bits_tag;
  wire [31:0] dcacheArb_io_requestor_1_resp_bits_data;
  wire  dcacheArb_io_requestor_1_resp_bits_replay;
  wire  dcacheArb_io_requestor_1_resp_bits_has_data;
  wire [31:0] dcacheArb_io_requestor_1_resp_bits_data_word_bypass;
  wire  dcacheArb_io_requestor_1_replay_next;
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  wire  dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  wire  dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_ld;
  wire  dcacheArb_io_requestor_1_s2_xcpt_ae_st;
  wire  dcacheArb_io_requestor_1_invalidate_lr;
  wire  dcacheArb_io_requestor_1_ordered;
  wire  dcacheArb_io_mem_req_ready;
  wire  dcacheArb_io_mem_req_valid;
  wire [31:0] dcacheArb_io_mem_req_bits_addr;
  wire [6:0] dcacheArb_io_mem_req_bits_tag;
  wire [4:0] dcacheArb_io_mem_req_bits_cmd;
  wire [2:0] dcacheArb_io_mem_req_bits_typ;
  wire  dcacheArb_io_mem_req_bits_phys;
  wire  dcacheArb_io_mem_s1_kill;
  wire [31:0] dcacheArb_io_mem_s1_data_data;
  wire [3:0] dcacheArb_io_mem_s1_data_mask;
  wire  dcacheArb_io_mem_s2_nack;
  wire  dcacheArb_io_mem_resp_valid;
  wire [6:0] dcacheArb_io_mem_resp_bits_tag;
  wire [31:0] dcacheArb_io_mem_resp_bits_data;
  wire  dcacheArb_io_mem_resp_bits_replay;
  wire  dcacheArb_io_mem_resp_bits_has_data;
  wire [31:0] dcacheArb_io_mem_resp_bits_data_word_bypass;
  wire [31:0] dcacheArb_io_mem_resp_bits_data_raw;
  wire  dcacheArb_io_mem_replay_next;
  wire  dcacheArb_io_mem_s2_xcpt_ma_ld;
  wire  dcacheArb_io_mem_s2_xcpt_ma_st;
  wire  dcacheArb_io_mem_s2_xcpt_pf_ld;
  wire  dcacheArb_io_mem_s2_xcpt_pf_st;
  wire  dcacheArb_io_mem_s2_xcpt_ae_ld;
  wire  dcacheArb_io_mem_s2_xcpt_ae_st;
  wire  dcacheArb_io_mem_invalidate_lr;
  wire  dcacheArb_io_mem_ordered;
  wire  ptw_clock;
  wire  ptw_reset;
  wire  ptw_io_requestor_0_req_valid;
  wire [19:0] ptw_io_requestor_0_req_bits_addr;
  wire  ptw_io_requestor_0_resp_valid;
  wire [1:0] ptw_io_requestor_0_status_dprv;
  wire [1:0] ptw_io_requestor_0_status_prv;
  wire  ptw_io_requestor_0_status_mxr;
  wire  ptw_io_requestor_0_status_sum;
  wire  ptw_io_requestor_0_pmp_0_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_0_cfg_a;
  wire  ptw_io_requestor_0_pmp_0_cfg_x;
  wire  ptw_io_requestor_0_pmp_0_cfg_w;
  wire  ptw_io_requestor_0_pmp_0_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_0_addr;
  wire [31:0] ptw_io_requestor_0_pmp_0_mask;
  wire  ptw_io_requestor_0_pmp_1_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_1_cfg_a;
  wire  ptw_io_requestor_0_pmp_1_cfg_x;
  wire  ptw_io_requestor_0_pmp_1_cfg_w;
  wire  ptw_io_requestor_0_pmp_1_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_1_addr;
  wire [31:0] ptw_io_requestor_0_pmp_1_mask;
  wire  ptw_io_requestor_0_pmp_2_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_2_cfg_a;
  wire  ptw_io_requestor_0_pmp_2_cfg_x;
  wire  ptw_io_requestor_0_pmp_2_cfg_w;
  wire  ptw_io_requestor_0_pmp_2_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_2_addr;
  wire [31:0] ptw_io_requestor_0_pmp_2_mask;
  wire  ptw_io_requestor_0_pmp_3_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_3_cfg_a;
  wire  ptw_io_requestor_0_pmp_3_cfg_x;
  wire  ptw_io_requestor_0_pmp_3_cfg_w;
  wire  ptw_io_requestor_0_pmp_3_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_3_addr;
  wire [31:0] ptw_io_requestor_0_pmp_3_mask;
  wire  ptw_io_requestor_0_pmp_4_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_4_cfg_a;
  wire  ptw_io_requestor_0_pmp_4_cfg_x;
  wire  ptw_io_requestor_0_pmp_4_cfg_w;
  wire  ptw_io_requestor_0_pmp_4_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_4_addr;
  wire [31:0] ptw_io_requestor_0_pmp_4_mask;
  wire  ptw_io_requestor_0_pmp_5_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_5_cfg_a;
  wire  ptw_io_requestor_0_pmp_5_cfg_x;
  wire  ptw_io_requestor_0_pmp_5_cfg_w;
  wire  ptw_io_requestor_0_pmp_5_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_5_addr;
  wire [31:0] ptw_io_requestor_0_pmp_5_mask;
  wire  ptw_io_requestor_0_pmp_6_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_6_cfg_a;
  wire  ptw_io_requestor_0_pmp_6_cfg_x;
  wire  ptw_io_requestor_0_pmp_6_cfg_w;
  wire  ptw_io_requestor_0_pmp_6_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_6_addr;
  wire [31:0] ptw_io_requestor_0_pmp_6_mask;
  wire  ptw_io_requestor_0_pmp_7_cfg_l;
  wire [1:0] ptw_io_requestor_0_pmp_7_cfg_a;
  wire  ptw_io_requestor_0_pmp_7_cfg_x;
  wire  ptw_io_requestor_0_pmp_7_cfg_w;
  wire  ptw_io_requestor_0_pmp_7_cfg_r;
  wire [29:0] ptw_io_requestor_0_pmp_7_addr;
  wire [31:0] ptw_io_requestor_0_pmp_7_mask;
  wire  ptw_io_requestor_1_req_valid;
  wire [19:0] ptw_io_requestor_1_req_bits_addr;
  wire  ptw_io_requestor_1_resp_valid;
  wire [1:0] ptw_io_requestor_1_status_dprv;
  wire [1:0] ptw_io_requestor_1_status_prv;
  wire  ptw_io_requestor_1_status_mxr;
  wire  ptw_io_requestor_1_status_sum;
  wire  ptw_io_requestor_1_pmp_0_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_0_cfg_a;
  wire  ptw_io_requestor_1_pmp_0_cfg_x;
  wire  ptw_io_requestor_1_pmp_0_cfg_w;
  wire  ptw_io_requestor_1_pmp_0_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_0_addr;
  wire [31:0] ptw_io_requestor_1_pmp_0_mask;
  wire  ptw_io_requestor_1_pmp_1_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_1_cfg_a;
  wire  ptw_io_requestor_1_pmp_1_cfg_x;
  wire  ptw_io_requestor_1_pmp_1_cfg_w;
  wire  ptw_io_requestor_1_pmp_1_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_1_addr;
  wire [31:0] ptw_io_requestor_1_pmp_1_mask;
  wire  ptw_io_requestor_1_pmp_2_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_2_cfg_a;
  wire  ptw_io_requestor_1_pmp_2_cfg_x;
  wire  ptw_io_requestor_1_pmp_2_cfg_w;
  wire  ptw_io_requestor_1_pmp_2_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_2_addr;
  wire [31:0] ptw_io_requestor_1_pmp_2_mask;
  wire  ptw_io_requestor_1_pmp_3_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_3_cfg_a;
  wire  ptw_io_requestor_1_pmp_3_cfg_x;
  wire  ptw_io_requestor_1_pmp_3_cfg_w;
  wire  ptw_io_requestor_1_pmp_3_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_3_addr;
  wire [31:0] ptw_io_requestor_1_pmp_3_mask;
  wire  ptw_io_requestor_1_pmp_4_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_4_cfg_a;
  wire  ptw_io_requestor_1_pmp_4_cfg_x;
  wire  ptw_io_requestor_1_pmp_4_cfg_w;
  wire  ptw_io_requestor_1_pmp_4_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_4_addr;
  wire [31:0] ptw_io_requestor_1_pmp_4_mask;
  wire  ptw_io_requestor_1_pmp_5_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_5_cfg_a;
  wire  ptw_io_requestor_1_pmp_5_cfg_x;
  wire  ptw_io_requestor_1_pmp_5_cfg_w;
  wire  ptw_io_requestor_1_pmp_5_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_5_addr;
  wire [31:0] ptw_io_requestor_1_pmp_5_mask;
  wire  ptw_io_requestor_1_pmp_6_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_6_cfg_a;
  wire  ptw_io_requestor_1_pmp_6_cfg_x;
  wire  ptw_io_requestor_1_pmp_6_cfg_w;
  wire  ptw_io_requestor_1_pmp_6_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_6_addr;
  wire [31:0] ptw_io_requestor_1_pmp_6_mask;
  wire  ptw_io_requestor_1_pmp_7_cfg_l;
  wire [1:0] ptw_io_requestor_1_pmp_7_cfg_a;
  wire  ptw_io_requestor_1_pmp_7_cfg_x;
  wire  ptw_io_requestor_1_pmp_7_cfg_w;
  wire  ptw_io_requestor_1_pmp_7_cfg_r;
  wire [29:0] ptw_io_requestor_1_pmp_7_addr;
  wire [31:0] ptw_io_requestor_1_pmp_7_mask;
  wire  ptw_io_mem_req_ready;
  wire  ptw_io_mem_s2_nack;
  wire  ptw_io_mem_resp_valid;
  wire [31:0] ptw_io_mem_resp_bits_data;
  wire  ptw_io_mem_s2_xcpt_ae_ld;
  wire [21:0] ptw_io_dpath_ptbr_ppn;
  wire  ptw_io_dpath_sfence_valid;
  wire  ptw_io_dpath_sfence_bits_rs1;
  wire [1:0] ptw_io_dpath_status_dprv;
  wire [1:0] ptw_io_dpath_status_prv;
  wire  ptw_io_dpath_status_mxr;
  wire  ptw_io_dpath_status_sum;
  wire  ptw_io_dpath_pmp_0_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_0_cfg_a;
  wire  ptw_io_dpath_pmp_0_cfg_x;
  wire  ptw_io_dpath_pmp_0_cfg_w;
  wire  ptw_io_dpath_pmp_0_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_0_addr;
  wire [31:0] ptw_io_dpath_pmp_0_mask;
  wire  ptw_io_dpath_pmp_1_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_1_cfg_a;
  wire  ptw_io_dpath_pmp_1_cfg_x;
  wire  ptw_io_dpath_pmp_1_cfg_w;
  wire  ptw_io_dpath_pmp_1_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_1_addr;
  wire [31:0] ptw_io_dpath_pmp_1_mask;
  wire  ptw_io_dpath_pmp_2_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_2_cfg_a;
  wire  ptw_io_dpath_pmp_2_cfg_x;
  wire  ptw_io_dpath_pmp_2_cfg_w;
  wire  ptw_io_dpath_pmp_2_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_2_addr;
  wire [31:0] ptw_io_dpath_pmp_2_mask;
  wire  ptw_io_dpath_pmp_3_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_3_cfg_a;
  wire  ptw_io_dpath_pmp_3_cfg_x;
  wire  ptw_io_dpath_pmp_3_cfg_w;
  wire  ptw_io_dpath_pmp_3_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_3_addr;
  wire [31:0] ptw_io_dpath_pmp_3_mask;
  wire  ptw_io_dpath_pmp_4_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_4_cfg_a;
  wire  ptw_io_dpath_pmp_4_cfg_x;
  wire  ptw_io_dpath_pmp_4_cfg_w;
  wire  ptw_io_dpath_pmp_4_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_4_addr;
  wire [31:0] ptw_io_dpath_pmp_4_mask;
  wire  ptw_io_dpath_pmp_5_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_5_cfg_a;
  wire  ptw_io_dpath_pmp_5_cfg_x;
  wire  ptw_io_dpath_pmp_5_cfg_w;
  wire  ptw_io_dpath_pmp_5_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_5_addr;
  wire [31:0] ptw_io_dpath_pmp_5_mask;
  wire  ptw_io_dpath_pmp_6_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_6_cfg_a;
  wire  ptw_io_dpath_pmp_6_cfg_x;
  wire  ptw_io_dpath_pmp_6_cfg_w;
  wire  ptw_io_dpath_pmp_6_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_6_addr;
  wire [31:0] ptw_io_dpath_pmp_6_mask;
  wire  ptw_io_dpath_pmp_7_cfg_l;
  wire [1:0] ptw_io_dpath_pmp_7_cfg_a;
  wire  ptw_io_dpath_pmp_7_cfg_x;
  wire  ptw_io_dpath_pmp_7_cfg_w;
  wire  ptw_io_dpath_pmp_7_cfg_r;
  wire [29:0] ptw_io_dpath_pmp_7_addr;
  wire [31:0] ptw_io_dpath_pmp_7_mask;
  wire  core_clock;
  wire  core_reset;
  wire  core_io_hartid;
  wire  core_io_interrupts_debug;
  wire  core_io_interrupts_mtip;
  wire  core_io_interrupts_msip;
  wire  core_io_interrupts_meip;
  wire  core_io_imem_req_valid;
  wire [31:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_req_bits_speculative;
  wire  core_io_imem_sfence_valid;
  wire  core_io_imem_sfence_bits_rs1;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire  core_io_imem_resp_bits_btb_valid;
  wire  core_io_imem_resp_bits_btb_bits_taken;
  wire  core_io_imem_resp_bits_btb_bits_bridx;
  wire [31:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data;
  wire  core_io_imem_resp_bits_xcpt_pf_inst;
  wire  core_io_imem_resp_bits_xcpt_ae_inst;
  wire  core_io_imem_resp_bits_replay;
  wire  core_io_imem_flush_icache;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [31:0] core_io_dmem_req_bits_addr;
  wire [6:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire  core_io_dmem_s1_kill;
  wire [31:0] core_io_dmem_s1_data_data;
  wire [3:0] core_io_dmem_s1_data_mask;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [6:0] core_io_dmem_resp_bits_tag;
  wire [31:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [31:0] core_io_dmem_resp_bits_data_word_bypass;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_s2_xcpt_ma_ld;
  wire  core_io_dmem_s2_xcpt_ma_st;
  wire  core_io_dmem_s2_xcpt_pf_ld;
  wire  core_io_dmem_s2_xcpt_pf_st;
  wire  core_io_dmem_s2_xcpt_ae_ld;
  wire  core_io_dmem_s2_xcpt_ae_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [21:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_sfence_valid;
  wire  core_io_ptw_sfence_bits_rs1;
  wire [1:0] core_io_ptw_status_dprv;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_mxr;
  wire  core_io_ptw_status_sum;
  wire  core_io_ptw_pmp_0_cfg_l;
  wire [1:0] core_io_ptw_pmp_0_cfg_a;
  wire  core_io_ptw_pmp_0_cfg_x;
  wire  core_io_ptw_pmp_0_cfg_w;
  wire  core_io_ptw_pmp_0_cfg_r;
  wire [29:0] core_io_ptw_pmp_0_addr;
  wire [31:0] core_io_ptw_pmp_0_mask;
  wire  core_io_ptw_pmp_1_cfg_l;
  wire [1:0] core_io_ptw_pmp_1_cfg_a;
  wire  core_io_ptw_pmp_1_cfg_x;
  wire  core_io_ptw_pmp_1_cfg_w;
  wire  core_io_ptw_pmp_1_cfg_r;
  wire [29:0] core_io_ptw_pmp_1_addr;
  wire [31:0] core_io_ptw_pmp_1_mask;
  wire  core_io_ptw_pmp_2_cfg_l;
  wire [1:0] core_io_ptw_pmp_2_cfg_a;
  wire  core_io_ptw_pmp_2_cfg_x;
  wire  core_io_ptw_pmp_2_cfg_w;
  wire  core_io_ptw_pmp_2_cfg_r;
  wire [29:0] core_io_ptw_pmp_2_addr;
  wire [31:0] core_io_ptw_pmp_2_mask;
  wire  core_io_ptw_pmp_3_cfg_l;
  wire [1:0] core_io_ptw_pmp_3_cfg_a;
  wire  core_io_ptw_pmp_3_cfg_x;
  wire  core_io_ptw_pmp_3_cfg_w;
  wire  core_io_ptw_pmp_3_cfg_r;
  wire [29:0] core_io_ptw_pmp_3_addr;
  wire [31:0] core_io_ptw_pmp_3_mask;
  wire  core_io_ptw_pmp_4_cfg_l;
  wire [1:0] core_io_ptw_pmp_4_cfg_a;
  wire  core_io_ptw_pmp_4_cfg_x;
  wire  core_io_ptw_pmp_4_cfg_w;
  wire  core_io_ptw_pmp_4_cfg_r;
  wire [29:0] core_io_ptw_pmp_4_addr;
  wire [31:0] core_io_ptw_pmp_4_mask;
  wire  core_io_ptw_pmp_5_cfg_l;
  wire [1:0] core_io_ptw_pmp_5_cfg_a;
  wire  core_io_ptw_pmp_5_cfg_x;
  wire  core_io_ptw_pmp_5_cfg_w;
  wire  core_io_ptw_pmp_5_cfg_r;
  wire [29:0] core_io_ptw_pmp_5_addr;
  wire [31:0] core_io_ptw_pmp_5_mask;
  wire  core_io_ptw_pmp_6_cfg_l;
  wire [1:0] core_io_ptw_pmp_6_cfg_a;
  wire  core_io_ptw_pmp_6_cfg_x;
  wire  core_io_ptw_pmp_6_cfg_w;
  wire  core_io_ptw_pmp_6_cfg_r;
  wire [29:0] core_io_ptw_pmp_6_addr;
  wire [31:0] core_io_ptw_pmp_6_mask;
  wire  core_io_ptw_pmp_7_cfg_l;
  wire [1:0] core_io_ptw_pmp_7_cfg_a;
  wire  core_io_ptw_pmp_7_cfg_x;
  wire  core_io_ptw_pmp_7_cfg_w;
  wire  core_io_ptw_pmp_7_cfg_r;
  wire [29:0] core_io_ptw_pmp_7_addr;
  wire [31:0] core_io_ptw_pmp_7_mask;
  wire [31:0] core_io_fpu_store_data;
  wire [31:0] core_io_fpu_toint_data;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_interrupt;
  TLXbar_tileBus tileBus (
    .clock(tileBus_clock),
    .reset(tileBus_reset),
    .io_in_1_a_ready(tileBus_io_in_1_a_ready),
    .io_in_1_a_valid(tileBus_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(tileBus_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_param(tileBus_io_in_1_a_bits_param),
    .io_in_1_a_bits_size(tileBus_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(tileBus_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(tileBus_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(tileBus_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(tileBus_io_in_1_a_bits_data),
    .io_in_1_d_ready(tileBus_io_in_1_d_ready),
    .io_in_1_d_valid(tileBus_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(tileBus_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_size(tileBus_io_in_1_d_bits_size),
    .io_in_1_d_bits_data(tileBus_io_in_1_d_bits_data),
    .io_in_1_d_bits_error(tileBus_io_in_1_d_bits_error),
    .io_in_0_a_ready(tileBus_io_in_0_a_ready),
    .io_in_0_a_valid(tileBus_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(tileBus_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(tileBus_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(tileBus_io_in_0_a_bits_size),
    .io_in_0_a_bits_address(tileBus_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(tileBus_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(tileBus_io_in_0_a_bits_data),
    .io_in_0_b_valid(tileBus_io_in_0_b_valid),
    .io_in_0_b_bits_param(tileBus_io_in_0_b_bits_param),
    .io_in_0_b_bits_address(tileBus_io_in_0_b_bits_address),
    .io_in_0_c_ready(tileBus_io_in_0_c_ready),
    .io_in_0_d_ready(tileBus_io_in_0_d_ready),
    .io_in_0_d_valid(tileBus_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(tileBus_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(tileBus_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(tileBus_io_in_0_d_bits_source),
    .io_in_0_d_bits_data(tileBus_io_in_0_d_bits_data),
    .io_in_0_e_ready(tileBus_io_in_0_e_ready),
    .io_out_0_a_ready(tileBus_io_out_0_a_ready),
    .io_out_0_a_valid(tileBus_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(tileBus_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(tileBus_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(tileBus_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(tileBus_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(tileBus_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(tileBus_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(tileBus_io_out_0_a_bits_data),
    .io_out_0_d_ready(tileBus_io_out_0_d_ready),
    .io_out_0_d_valid(tileBus_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(tileBus_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(tileBus_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(tileBus_io_out_0_d_bits_source),
    .io_out_0_d_bits_data(tileBus_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(tileBus_io_out_0_d_bits_error)
  );
  DCache_dcache dcache (
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_cpu_req_ready(dcache_io_cpu_req_ready),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(dcache_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(dcache_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(dcache_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(dcache_io_cpu_req_bits_phys),
    .io_cpu_s1_kill(dcache_io_cpu_s1_kill),
    .io_cpu_s1_data_data(dcache_io_cpu_s1_data_data),
    .io_cpu_s1_data_mask(dcache_io_cpu_s1_data_mask),
    .io_cpu_s2_nack(dcache_io_cpu_s2_nack),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_tag(dcache_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(dcache_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(dcache_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(dcache_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_data_raw(dcache_io_cpu_resp_bits_data_raw),
    .io_cpu_replay_next(dcache_io_cpu_replay_next),
    .io_cpu_s2_xcpt_ma_ld(dcache_io_cpu_s2_xcpt_ma_ld),
    .io_cpu_s2_xcpt_ma_st(dcache_io_cpu_s2_xcpt_ma_st),
    .io_cpu_s2_xcpt_pf_ld(dcache_io_cpu_s2_xcpt_pf_ld),
    .io_cpu_s2_xcpt_pf_st(dcache_io_cpu_s2_xcpt_pf_st),
    .io_cpu_s2_xcpt_ae_ld(dcache_io_cpu_s2_xcpt_ae_ld),
    .io_cpu_s2_xcpt_ae_st(dcache_io_cpu_s2_xcpt_ae_st),
    .io_cpu_invalidate_lr(dcache_io_cpu_invalidate_lr),
    .io_cpu_ordered(dcache_io_cpu_ordered),
    .io_ptw_req_valid(dcache_io_ptw_req_valid),
    .io_ptw_req_bits_addr(dcache_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(dcache_io_ptw_resp_valid),
    .io_ptw_status_dprv(dcache_io_ptw_status_dprv),
    .io_ptw_status_prv(dcache_io_ptw_status_prv),
    .io_ptw_status_mxr(dcache_io_ptw_status_mxr),
    .io_ptw_status_sum(dcache_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(dcache_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(dcache_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(dcache_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(dcache_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(dcache_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(dcache_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(dcache_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(dcache_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(dcache_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(dcache_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(dcache_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(dcache_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(dcache_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(dcache_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(dcache_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(dcache_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(dcache_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(dcache_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(dcache_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(dcache_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(dcache_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(dcache_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(dcache_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(dcache_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(dcache_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(dcache_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(dcache_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(dcache_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(dcache_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(dcache_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(dcache_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(dcache_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(dcache_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(dcache_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(dcache_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(dcache_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(dcache_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(dcache_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(dcache_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(dcache_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(dcache_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(dcache_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(dcache_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(dcache_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(dcache_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(dcache_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(dcache_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(dcache_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(dcache_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(dcache_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(dcache_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(dcache_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(dcache_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(dcache_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(dcache_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(dcache_io_ptw_pmp_7_mask),
    .io_mem_0_a_ready(dcache_io_mem_0_a_ready),
    .io_mem_0_a_valid(dcache_io_mem_0_a_valid),
    .io_mem_0_a_bits_opcode(dcache_io_mem_0_a_bits_opcode),
    .io_mem_0_a_bits_param(dcache_io_mem_0_a_bits_param),
    .io_mem_0_a_bits_size(dcache_io_mem_0_a_bits_size),
    .io_mem_0_a_bits_address(dcache_io_mem_0_a_bits_address),
    .io_mem_0_a_bits_mask(dcache_io_mem_0_a_bits_mask),
    .io_mem_0_a_bits_data(dcache_io_mem_0_a_bits_data),
    .io_mem_0_b_ready(dcache_io_mem_0_b_ready),
    .io_mem_0_b_valid(dcache_io_mem_0_b_valid),
    .io_mem_0_b_bits_param(dcache_io_mem_0_b_bits_param),
    .io_mem_0_b_bits_address(dcache_io_mem_0_b_bits_address),
    .io_mem_0_c_ready(dcache_io_mem_0_c_ready),
    .io_mem_0_c_valid(dcache_io_mem_0_c_valid),
    .io_mem_0_c_bits_address(dcache_io_mem_0_c_bits_address),
    .io_mem_0_d_ready(dcache_io_mem_0_d_ready),
    .io_mem_0_d_valid(dcache_io_mem_0_d_valid),
    .io_mem_0_d_bits_opcode(dcache_io_mem_0_d_bits_opcode),
    .io_mem_0_d_bits_size(dcache_io_mem_0_d_bits_size),
    .io_mem_0_d_bits_source(dcache_io_mem_0_d_bits_source),
    .io_mem_0_d_bits_data(dcache_io_mem_0_d_bits_data),
    .io_mem_0_e_ready(dcache_io_mem_0_e_ready),
    .io_mem_0_e_valid(dcache_io_mem_0_e_valid)
  );
  Frontend_frontend frontend (
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_tl_out_0_a_ready(frontend_io_tl_out_0_a_ready),
    .io_tl_out_0_a_valid(frontend_io_tl_out_0_a_valid),
    .io_tl_out_0_a_bits_opcode(frontend_io_tl_out_0_a_bits_opcode),
    .io_tl_out_0_a_bits_param(frontend_io_tl_out_0_a_bits_param),
    .io_tl_out_0_a_bits_size(frontend_io_tl_out_0_a_bits_size),
    .io_tl_out_0_a_bits_source(frontend_io_tl_out_0_a_bits_source),
    .io_tl_out_0_a_bits_address(frontend_io_tl_out_0_a_bits_address),
    .io_tl_out_0_a_bits_mask(frontend_io_tl_out_0_a_bits_mask),
    .io_tl_out_0_a_bits_data(frontend_io_tl_out_0_a_bits_data),
    .io_tl_out_0_d_ready(frontend_io_tl_out_0_d_ready),
    .io_tl_out_0_d_valid(frontend_io_tl_out_0_d_valid),
    .io_tl_out_0_d_bits_opcode(frontend_io_tl_out_0_d_bits_opcode),
    .io_tl_out_0_d_bits_size(frontend_io_tl_out_0_d_bits_size),
    .io_tl_out_0_d_bits_data(frontend_io_tl_out_0_d_bits_data),
    .io_tl_out_0_d_bits_error(frontend_io_tl_out_0_d_bits_error),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(frontend_io_cpu_req_bits_speculative),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_btb_valid(frontend_io_cpu_resp_bits_btb_valid),
    .io_cpu_resp_bits_btb_bits_taken(frontend_io_cpu_resp_bits_btb_bits_taken),
    .io_cpu_resp_bits_btb_bits_bridx(frontend_io_cpu_resp_bits_btb_bits_bridx),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data(frontend_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_xcpt_pf_inst(frontend_io_cpu_resp_bits_xcpt_pf_inst),
    .io_cpu_resp_bits_xcpt_ae_inst(frontend_io_cpu_resp_bits_xcpt_ae_inst),
    .io_cpu_resp_bits_replay(frontend_io_cpu_resp_bits_replay),
    .io_cpu_flush_icache(frontend_io_cpu_flush_icache),
    .io_cpu_npc(frontend_io_cpu_npc),
    .io_ptw_req_valid(frontend_io_ptw_req_valid),
    .io_ptw_req_bits_addr(frontend_io_ptw_req_bits_addr),
    .io_ptw_resp_valid(frontend_io_ptw_resp_valid),
    .io_ptw_status_dprv(frontend_io_ptw_status_dprv),
    .io_ptw_status_prv(frontend_io_ptw_status_prv),
    .io_ptw_status_mxr(frontend_io_ptw_status_mxr),
    .io_ptw_status_sum(frontend_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(frontend_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(frontend_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(frontend_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(frontend_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(frontend_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(frontend_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(frontend_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(frontend_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(frontend_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(frontend_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(frontend_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(frontend_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(frontend_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(frontend_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(frontend_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(frontend_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(frontend_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(frontend_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(frontend_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(frontend_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(frontend_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(frontend_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(frontend_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(frontend_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(frontend_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(frontend_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(frontend_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(frontend_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(frontend_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(frontend_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(frontend_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(frontend_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(frontend_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(frontend_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(frontend_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(frontend_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(frontend_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(frontend_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(frontend_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(frontend_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(frontend_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(frontend_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(frontend_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(frontend_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(frontend_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(frontend_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(frontend_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(frontend_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(frontend_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(frontend_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(frontend_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(frontend_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(frontend_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(frontend_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(frontend_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(frontend_io_ptw_pmp_7_mask),
    .io_resetVector(frontend_io_resetVector)
  );
  ScratchpadSlavePort ScratchpadSlavePort (
    .clock(ScratchpadSlavePort_clock),
    .reset(ScratchpadSlavePort_reset),
    .io_tl_in_0_a_ready(ScratchpadSlavePort_io_tl_in_0_a_ready),
    .io_tl_in_0_a_valid(ScratchpadSlavePort_io_tl_in_0_a_valid),
    .io_tl_in_0_a_bits_opcode(ScratchpadSlavePort_io_tl_in_0_a_bits_opcode),
    .io_tl_in_0_a_bits_param(ScratchpadSlavePort_io_tl_in_0_a_bits_param),
    .io_tl_in_0_a_bits_size(ScratchpadSlavePort_io_tl_in_0_a_bits_size),
    .io_tl_in_0_a_bits_source(ScratchpadSlavePort_io_tl_in_0_a_bits_source),
    .io_tl_in_0_a_bits_address(ScratchpadSlavePort_io_tl_in_0_a_bits_address),
    .io_tl_in_0_a_bits_mask(ScratchpadSlavePort_io_tl_in_0_a_bits_mask),
    .io_tl_in_0_a_bits_data(ScratchpadSlavePort_io_tl_in_0_a_bits_data),
    .io_tl_in_0_d_ready(ScratchpadSlavePort_io_tl_in_0_d_ready),
    .io_tl_in_0_d_valid(ScratchpadSlavePort_io_tl_in_0_d_valid),
    .io_tl_in_0_d_bits_opcode(ScratchpadSlavePort_io_tl_in_0_d_bits_opcode),
    .io_tl_in_0_d_bits_param(ScratchpadSlavePort_io_tl_in_0_d_bits_param),
    .io_tl_in_0_d_bits_size(ScratchpadSlavePort_io_tl_in_0_d_bits_size),
    .io_tl_in_0_d_bits_source(ScratchpadSlavePort_io_tl_in_0_d_bits_source),
    .io_tl_in_0_d_bits_sink(ScratchpadSlavePort_io_tl_in_0_d_bits_sink),
    .io_tl_in_0_d_bits_data(ScratchpadSlavePort_io_tl_in_0_d_bits_data),
    .io_tl_in_0_d_bits_error(ScratchpadSlavePort_io_tl_in_0_d_bits_error),
    .io_dmem_req_ready(ScratchpadSlavePort_io_dmem_req_ready),
    .io_dmem_req_valid(ScratchpadSlavePort_io_dmem_req_valid),
    .io_dmem_req_bits_addr(ScratchpadSlavePort_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(ScratchpadSlavePort_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(ScratchpadSlavePort_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(ScratchpadSlavePort_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(ScratchpadSlavePort_io_dmem_req_bits_phys),
    .io_dmem_s1_kill(ScratchpadSlavePort_io_dmem_s1_kill),
    .io_dmem_s1_data_data(ScratchpadSlavePort_io_dmem_s1_data_data),
    .io_dmem_s1_data_mask(ScratchpadSlavePort_io_dmem_s1_data_mask),
    .io_dmem_s2_nack(ScratchpadSlavePort_io_dmem_s2_nack),
    .io_dmem_resp_valid(ScratchpadSlavePort_io_dmem_resp_valid),
    .io_dmem_resp_bits_data_raw(ScratchpadSlavePort_io_dmem_resp_bits_data_raw),
    .io_dmem_invalidate_lr(ScratchpadSlavePort_io_dmem_invalidate_lr)
  );
  TLFragmenter_2 TLFragmenter (
    .clock(TLFragmenter_clock),
    .reset(TLFragmenter_reset),
    .io_in_0_a_ready(TLFragmenter_io_in_0_a_ready),
    .io_in_0_a_valid(TLFragmenter_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLFragmenter_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLFragmenter_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLFragmenter_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLFragmenter_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLFragmenter_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLFragmenter_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLFragmenter_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLFragmenter_io_in_0_d_ready),
    .io_in_0_d_valid(TLFragmenter_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLFragmenter_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLFragmenter_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLFragmenter_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLFragmenter_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLFragmenter_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLFragmenter_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLFragmenter_io_in_0_d_bits_error),
    .io_out_0_a_ready(TLFragmenter_io_out_0_a_ready),
    .io_out_0_a_valid(TLFragmenter_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLFragmenter_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLFragmenter_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLFragmenter_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLFragmenter_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLFragmenter_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLFragmenter_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLFragmenter_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLFragmenter_io_out_0_d_ready),
    .io_out_0_d_valid(TLFragmenter_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLFragmenter_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLFragmenter_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLFragmenter_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLFragmenter_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLFragmenter_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLFragmenter_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLFragmenter_io_out_0_d_bits_error)
  );
  HellaCacheArbiter dcacheArb (
    .clock(dcacheArb_clock),
    .io_requestor_0_req_ready(dcacheArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcacheArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcacheArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcacheArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcacheArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcacheArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcacheArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_s1_kill(dcacheArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data_data(dcacheArb_io_requestor_0_s1_data_data),
    .io_requestor_0_s1_data_mask(dcacheArb_io_requestor_0_s1_data_mask),
    .io_requestor_0_s2_nack(dcacheArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcacheArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_data_raw(dcacheArb_io_requestor_0_resp_bits_data_raw),
    .io_requestor_0_invalidate_lr(dcacheArb_io_requestor_0_invalidate_lr),
    .io_requestor_1_req_ready(dcacheArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcacheArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcacheArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcacheArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcacheArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_typ(dcacheArb_io_requestor_1_req_bits_typ),
    .io_requestor_1_req_bits_phys(dcacheArb_io_requestor_1_req_bits_phys),
    .io_requestor_1_s1_kill(dcacheArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data_data(dcacheArb_io_requestor_1_s1_data_data),
    .io_requestor_1_s1_data_mask(dcacheArb_io_requestor_1_s1_data_mask),
    .io_requestor_1_s2_nack(dcacheArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcacheArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_tag(dcacheArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_data(dcacheArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcacheArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcacheArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcacheArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_replay_next(dcacheArb_io_requestor_1_replay_next),
    .io_requestor_1_s2_xcpt_ma_ld(dcacheArb_io_requestor_1_s2_xcpt_ma_ld),
    .io_requestor_1_s2_xcpt_ma_st(dcacheArb_io_requestor_1_s2_xcpt_ma_st),
    .io_requestor_1_s2_xcpt_pf_ld(dcacheArb_io_requestor_1_s2_xcpt_pf_ld),
    .io_requestor_1_s2_xcpt_pf_st(dcacheArb_io_requestor_1_s2_xcpt_pf_st),
    .io_requestor_1_s2_xcpt_ae_ld(dcacheArb_io_requestor_1_s2_xcpt_ae_ld),
    .io_requestor_1_s2_xcpt_ae_st(dcacheArb_io_requestor_1_s2_xcpt_ae_st),
    .io_requestor_1_invalidate_lr(dcacheArb_io_requestor_1_invalidate_lr),
    .io_requestor_1_ordered(dcacheArb_io_requestor_1_ordered),
    .io_mem_req_ready(dcacheArb_io_mem_req_ready),
    .io_mem_req_valid(dcacheArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcacheArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcacheArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcacheArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcacheArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcacheArb_io_mem_req_bits_phys),
    .io_mem_s1_kill(dcacheArb_io_mem_s1_kill),
    .io_mem_s1_data_data(dcacheArb_io_mem_s1_data_data),
    .io_mem_s1_data_mask(dcacheArb_io_mem_s1_data_mask),
    .io_mem_s2_nack(dcacheArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcacheArb_io_mem_resp_valid),
    .io_mem_resp_bits_tag(dcacheArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_data(dcacheArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcacheArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcacheArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcacheArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_data_raw(dcacheArb_io_mem_resp_bits_data_raw),
    .io_mem_replay_next(dcacheArb_io_mem_replay_next),
    .io_mem_s2_xcpt_ma_ld(dcacheArb_io_mem_s2_xcpt_ma_ld),
    .io_mem_s2_xcpt_ma_st(dcacheArb_io_mem_s2_xcpt_ma_st),
    .io_mem_s2_xcpt_pf_ld(dcacheArb_io_mem_s2_xcpt_pf_ld),
    .io_mem_s2_xcpt_pf_st(dcacheArb_io_mem_s2_xcpt_pf_st),
    .io_mem_s2_xcpt_ae_ld(dcacheArb_io_mem_s2_xcpt_ae_ld),
    .io_mem_s2_xcpt_ae_st(dcacheArb_io_mem_s2_xcpt_ae_st),
    .io_mem_invalidate_lr(dcacheArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcacheArb_io_mem_ordered)
  );
  PTW ptw (
    .clock(ptw_clock),
    .reset(ptw_reset),
    .io_requestor_0_req_valid(ptw_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(ptw_io_requestor_0_req_bits_addr),
    .io_requestor_0_resp_valid(ptw_io_requestor_0_resp_valid),
    .io_requestor_0_status_dprv(ptw_io_requestor_0_status_dprv),
    .io_requestor_0_status_prv(ptw_io_requestor_0_status_prv),
    .io_requestor_0_status_mxr(ptw_io_requestor_0_status_mxr),
    .io_requestor_0_status_sum(ptw_io_requestor_0_status_sum),
    .io_requestor_0_pmp_0_cfg_l(ptw_io_requestor_0_pmp_0_cfg_l),
    .io_requestor_0_pmp_0_cfg_a(ptw_io_requestor_0_pmp_0_cfg_a),
    .io_requestor_0_pmp_0_cfg_x(ptw_io_requestor_0_pmp_0_cfg_x),
    .io_requestor_0_pmp_0_cfg_w(ptw_io_requestor_0_pmp_0_cfg_w),
    .io_requestor_0_pmp_0_cfg_r(ptw_io_requestor_0_pmp_0_cfg_r),
    .io_requestor_0_pmp_0_addr(ptw_io_requestor_0_pmp_0_addr),
    .io_requestor_0_pmp_0_mask(ptw_io_requestor_0_pmp_0_mask),
    .io_requestor_0_pmp_1_cfg_l(ptw_io_requestor_0_pmp_1_cfg_l),
    .io_requestor_0_pmp_1_cfg_a(ptw_io_requestor_0_pmp_1_cfg_a),
    .io_requestor_0_pmp_1_cfg_x(ptw_io_requestor_0_pmp_1_cfg_x),
    .io_requestor_0_pmp_1_cfg_w(ptw_io_requestor_0_pmp_1_cfg_w),
    .io_requestor_0_pmp_1_cfg_r(ptw_io_requestor_0_pmp_1_cfg_r),
    .io_requestor_0_pmp_1_addr(ptw_io_requestor_0_pmp_1_addr),
    .io_requestor_0_pmp_1_mask(ptw_io_requestor_0_pmp_1_mask),
    .io_requestor_0_pmp_2_cfg_l(ptw_io_requestor_0_pmp_2_cfg_l),
    .io_requestor_0_pmp_2_cfg_a(ptw_io_requestor_0_pmp_2_cfg_a),
    .io_requestor_0_pmp_2_cfg_x(ptw_io_requestor_0_pmp_2_cfg_x),
    .io_requestor_0_pmp_2_cfg_w(ptw_io_requestor_0_pmp_2_cfg_w),
    .io_requestor_0_pmp_2_cfg_r(ptw_io_requestor_0_pmp_2_cfg_r),
    .io_requestor_0_pmp_2_addr(ptw_io_requestor_0_pmp_2_addr),
    .io_requestor_0_pmp_2_mask(ptw_io_requestor_0_pmp_2_mask),
    .io_requestor_0_pmp_3_cfg_l(ptw_io_requestor_0_pmp_3_cfg_l),
    .io_requestor_0_pmp_3_cfg_a(ptw_io_requestor_0_pmp_3_cfg_a),
    .io_requestor_0_pmp_3_cfg_x(ptw_io_requestor_0_pmp_3_cfg_x),
    .io_requestor_0_pmp_3_cfg_w(ptw_io_requestor_0_pmp_3_cfg_w),
    .io_requestor_0_pmp_3_cfg_r(ptw_io_requestor_0_pmp_3_cfg_r),
    .io_requestor_0_pmp_3_addr(ptw_io_requestor_0_pmp_3_addr),
    .io_requestor_0_pmp_3_mask(ptw_io_requestor_0_pmp_3_mask),
    .io_requestor_0_pmp_4_cfg_l(ptw_io_requestor_0_pmp_4_cfg_l),
    .io_requestor_0_pmp_4_cfg_a(ptw_io_requestor_0_pmp_4_cfg_a),
    .io_requestor_0_pmp_4_cfg_x(ptw_io_requestor_0_pmp_4_cfg_x),
    .io_requestor_0_pmp_4_cfg_w(ptw_io_requestor_0_pmp_4_cfg_w),
    .io_requestor_0_pmp_4_cfg_r(ptw_io_requestor_0_pmp_4_cfg_r),
    .io_requestor_0_pmp_4_addr(ptw_io_requestor_0_pmp_4_addr),
    .io_requestor_0_pmp_4_mask(ptw_io_requestor_0_pmp_4_mask),
    .io_requestor_0_pmp_5_cfg_l(ptw_io_requestor_0_pmp_5_cfg_l),
    .io_requestor_0_pmp_5_cfg_a(ptw_io_requestor_0_pmp_5_cfg_a),
    .io_requestor_0_pmp_5_cfg_x(ptw_io_requestor_0_pmp_5_cfg_x),
    .io_requestor_0_pmp_5_cfg_w(ptw_io_requestor_0_pmp_5_cfg_w),
    .io_requestor_0_pmp_5_cfg_r(ptw_io_requestor_0_pmp_5_cfg_r),
    .io_requestor_0_pmp_5_addr(ptw_io_requestor_0_pmp_5_addr),
    .io_requestor_0_pmp_5_mask(ptw_io_requestor_0_pmp_5_mask),
    .io_requestor_0_pmp_6_cfg_l(ptw_io_requestor_0_pmp_6_cfg_l),
    .io_requestor_0_pmp_6_cfg_a(ptw_io_requestor_0_pmp_6_cfg_a),
    .io_requestor_0_pmp_6_cfg_x(ptw_io_requestor_0_pmp_6_cfg_x),
    .io_requestor_0_pmp_6_cfg_w(ptw_io_requestor_0_pmp_6_cfg_w),
    .io_requestor_0_pmp_6_cfg_r(ptw_io_requestor_0_pmp_6_cfg_r),
    .io_requestor_0_pmp_6_addr(ptw_io_requestor_0_pmp_6_addr),
    .io_requestor_0_pmp_6_mask(ptw_io_requestor_0_pmp_6_mask),
    .io_requestor_0_pmp_7_cfg_l(ptw_io_requestor_0_pmp_7_cfg_l),
    .io_requestor_0_pmp_7_cfg_a(ptw_io_requestor_0_pmp_7_cfg_a),
    .io_requestor_0_pmp_7_cfg_x(ptw_io_requestor_0_pmp_7_cfg_x),
    .io_requestor_0_pmp_7_cfg_w(ptw_io_requestor_0_pmp_7_cfg_w),
    .io_requestor_0_pmp_7_cfg_r(ptw_io_requestor_0_pmp_7_cfg_r),
    .io_requestor_0_pmp_7_addr(ptw_io_requestor_0_pmp_7_addr),
    .io_requestor_0_pmp_7_mask(ptw_io_requestor_0_pmp_7_mask),
    .io_requestor_1_req_valid(ptw_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(ptw_io_requestor_1_req_bits_addr),
    .io_requestor_1_resp_valid(ptw_io_requestor_1_resp_valid),
    .io_requestor_1_status_dprv(ptw_io_requestor_1_status_dprv),
    .io_requestor_1_status_prv(ptw_io_requestor_1_status_prv),
    .io_requestor_1_status_mxr(ptw_io_requestor_1_status_mxr),
    .io_requestor_1_status_sum(ptw_io_requestor_1_status_sum),
    .io_requestor_1_pmp_0_cfg_l(ptw_io_requestor_1_pmp_0_cfg_l),
    .io_requestor_1_pmp_0_cfg_a(ptw_io_requestor_1_pmp_0_cfg_a),
    .io_requestor_1_pmp_0_cfg_x(ptw_io_requestor_1_pmp_0_cfg_x),
    .io_requestor_1_pmp_0_cfg_w(ptw_io_requestor_1_pmp_0_cfg_w),
    .io_requestor_1_pmp_0_cfg_r(ptw_io_requestor_1_pmp_0_cfg_r),
    .io_requestor_1_pmp_0_addr(ptw_io_requestor_1_pmp_0_addr),
    .io_requestor_1_pmp_0_mask(ptw_io_requestor_1_pmp_0_mask),
    .io_requestor_1_pmp_1_cfg_l(ptw_io_requestor_1_pmp_1_cfg_l),
    .io_requestor_1_pmp_1_cfg_a(ptw_io_requestor_1_pmp_1_cfg_a),
    .io_requestor_1_pmp_1_cfg_x(ptw_io_requestor_1_pmp_1_cfg_x),
    .io_requestor_1_pmp_1_cfg_w(ptw_io_requestor_1_pmp_1_cfg_w),
    .io_requestor_1_pmp_1_cfg_r(ptw_io_requestor_1_pmp_1_cfg_r),
    .io_requestor_1_pmp_1_addr(ptw_io_requestor_1_pmp_1_addr),
    .io_requestor_1_pmp_1_mask(ptw_io_requestor_1_pmp_1_mask),
    .io_requestor_1_pmp_2_cfg_l(ptw_io_requestor_1_pmp_2_cfg_l),
    .io_requestor_1_pmp_2_cfg_a(ptw_io_requestor_1_pmp_2_cfg_a),
    .io_requestor_1_pmp_2_cfg_x(ptw_io_requestor_1_pmp_2_cfg_x),
    .io_requestor_1_pmp_2_cfg_w(ptw_io_requestor_1_pmp_2_cfg_w),
    .io_requestor_1_pmp_2_cfg_r(ptw_io_requestor_1_pmp_2_cfg_r),
    .io_requestor_1_pmp_2_addr(ptw_io_requestor_1_pmp_2_addr),
    .io_requestor_1_pmp_2_mask(ptw_io_requestor_1_pmp_2_mask),
    .io_requestor_1_pmp_3_cfg_l(ptw_io_requestor_1_pmp_3_cfg_l),
    .io_requestor_1_pmp_3_cfg_a(ptw_io_requestor_1_pmp_3_cfg_a),
    .io_requestor_1_pmp_3_cfg_x(ptw_io_requestor_1_pmp_3_cfg_x),
    .io_requestor_1_pmp_3_cfg_w(ptw_io_requestor_1_pmp_3_cfg_w),
    .io_requestor_1_pmp_3_cfg_r(ptw_io_requestor_1_pmp_3_cfg_r),
    .io_requestor_1_pmp_3_addr(ptw_io_requestor_1_pmp_3_addr),
    .io_requestor_1_pmp_3_mask(ptw_io_requestor_1_pmp_3_mask),
    .io_requestor_1_pmp_4_cfg_l(ptw_io_requestor_1_pmp_4_cfg_l),
    .io_requestor_1_pmp_4_cfg_a(ptw_io_requestor_1_pmp_4_cfg_a),
    .io_requestor_1_pmp_4_cfg_x(ptw_io_requestor_1_pmp_4_cfg_x),
    .io_requestor_1_pmp_4_cfg_w(ptw_io_requestor_1_pmp_4_cfg_w),
    .io_requestor_1_pmp_4_cfg_r(ptw_io_requestor_1_pmp_4_cfg_r),
    .io_requestor_1_pmp_4_addr(ptw_io_requestor_1_pmp_4_addr),
    .io_requestor_1_pmp_4_mask(ptw_io_requestor_1_pmp_4_mask),
    .io_requestor_1_pmp_5_cfg_l(ptw_io_requestor_1_pmp_5_cfg_l),
    .io_requestor_1_pmp_5_cfg_a(ptw_io_requestor_1_pmp_5_cfg_a),
    .io_requestor_1_pmp_5_cfg_x(ptw_io_requestor_1_pmp_5_cfg_x),
    .io_requestor_1_pmp_5_cfg_w(ptw_io_requestor_1_pmp_5_cfg_w),
    .io_requestor_1_pmp_5_cfg_r(ptw_io_requestor_1_pmp_5_cfg_r),
    .io_requestor_1_pmp_5_addr(ptw_io_requestor_1_pmp_5_addr),
    .io_requestor_1_pmp_5_mask(ptw_io_requestor_1_pmp_5_mask),
    .io_requestor_1_pmp_6_cfg_l(ptw_io_requestor_1_pmp_6_cfg_l),
    .io_requestor_1_pmp_6_cfg_a(ptw_io_requestor_1_pmp_6_cfg_a),
    .io_requestor_1_pmp_6_cfg_x(ptw_io_requestor_1_pmp_6_cfg_x),
    .io_requestor_1_pmp_6_cfg_w(ptw_io_requestor_1_pmp_6_cfg_w),
    .io_requestor_1_pmp_6_cfg_r(ptw_io_requestor_1_pmp_6_cfg_r),
    .io_requestor_1_pmp_6_addr(ptw_io_requestor_1_pmp_6_addr),
    .io_requestor_1_pmp_6_mask(ptw_io_requestor_1_pmp_6_mask),
    .io_requestor_1_pmp_7_cfg_l(ptw_io_requestor_1_pmp_7_cfg_l),
    .io_requestor_1_pmp_7_cfg_a(ptw_io_requestor_1_pmp_7_cfg_a),
    .io_requestor_1_pmp_7_cfg_x(ptw_io_requestor_1_pmp_7_cfg_x),
    .io_requestor_1_pmp_7_cfg_w(ptw_io_requestor_1_pmp_7_cfg_w),
    .io_requestor_1_pmp_7_cfg_r(ptw_io_requestor_1_pmp_7_cfg_r),
    .io_requestor_1_pmp_7_addr(ptw_io_requestor_1_pmp_7_addr),
    .io_requestor_1_pmp_7_mask(ptw_io_requestor_1_pmp_7_mask),
    .io_mem_req_ready(ptw_io_mem_req_ready),
    .io_mem_s2_nack(ptw_io_mem_s2_nack),
    .io_mem_resp_valid(ptw_io_mem_resp_valid),
    .io_mem_resp_bits_data(ptw_io_mem_resp_bits_data),
    .io_mem_s2_xcpt_ae_ld(ptw_io_mem_s2_xcpt_ae_ld),
    .io_dpath_ptbr_ppn(ptw_io_dpath_ptbr_ppn),
    .io_dpath_sfence_valid(ptw_io_dpath_sfence_valid),
    .io_dpath_sfence_bits_rs1(ptw_io_dpath_sfence_bits_rs1),
    .io_dpath_status_dprv(ptw_io_dpath_status_dprv),
    .io_dpath_status_prv(ptw_io_dpath_status_prv),
    .io_dpath_status_mxr(ptw_io_dpath_status_mxr),
    .io_dpath_status_sum(ptw_io_dpath_status_sum),
    .io_dpath_pmp_0_cfg_l(ptw_io_dpath_pmp_0_cfg_l),
    .io_dpath_pmp_0_cfg_a(ptw_io_dpath_pmp_0_cfg_a),
    .io_dpath_pmp_0_cfg_x(ptw_io_dpath_pmp_0_cfg_x),
    .io_dpath_pmp_0_cfg_w(ptw_io_dpath_pmp_0_cfg_w),
    .io_dpath_pmp_0_cfg_r(ptw_io_dpath_pmp_0_cfg_r),
    .io_dpath_pmp_0_addr(ptw_io_dpath_pmp_0_addr),
    .io_dpath_pmp_0_mask(ptw_io_dpath_pmp_0_mask),
    .io_dpath_pmp_1_cfg_l(ptw_io_dpath_pmp_1_cfg_l),
    .io_dpath_pmp_1_cfg_a(ptw_io_dpath_pmp_1_cfg_a),
    .io_dpath_pmp_1_cfg_x(ptw_io_dpath_pmp_1_cfg_x),
    .io_dpath_pmp_1_cfg_w(ptw_io_dpath_pmp_1_cfg_w),
    .io_dpath_pmp_1_cfg_r(ptw_io_dpath_pmp_1_cfg_r),
    .io_dpath_pmp_1_addr(ptw_io_dpath_pmp_1_addr),
    .io_dpath_pmp_1_mask(ptw_io_dpath_pmp_1_mask),
    .io_dpath_pmp_2_cfg_l(ptw_io_dpath_pmp_2_cfg_l),
    .io_dpath_pmp_2_cfg_a(ptw_io_dpath_pmp_2_cfg_a),
    .io_dpath_pmp_2_cfg_x(ptw_io_dpath_pmp_2_cfg_x),
    .io_dpath_pmp_2_cfg_w(ptw_io_dpath_pmp_2_cfg_w),
    .io_dpath_pmp_2_cfg_r(ptw_io_dpath_pmp_2_cfg_r),
    .io_dpath_pmp_2_addr(ptw_io_dpath_pmp_2_addr),
    .io_dpath_pmp_2_mask(ptw_io_dpath_pmp_2_mask),
    .io_dpath_pmp_3_cfg_l(ptw_io_dpath_pmp_3_cfg_l),
    .io_dpath_pmp_3_cfg_a(ptw_io_dpath_pmp_3_cfg_a),
    .io_dpath_pmp_3_cfg_x(ptw_io_dpath_pmp_3_cfg_x),
    .io_dpath_pmp_3_cfg_w(ptw_io_dpath_pmp_3_cfg_w),
    .io_dpath_pmp_3_cfg_r(ptw_io_dpath_pmp_3_cfg_r),
    .io_dpath_pmp_3_addr(ptw_io_dpath_pmp_3_addr),
    .io_dpath_pmp_3_mask(ptw_io_dpath_pmp_3_mask),
    .io_dpath_pmp_4_cfg_l(ptw_io_dpath_pmp_4_cfg_l),
    .io_dpath_pmp_4_cfg_a(ptw_io_dpath_pmp_4_cfg_a),
    .io_dpath_pmp_4_cfg_x(ptw_io_dpath_pmp_4_cfg_x),
    .io_dpath_pmp_4_cfg_w(ptw_io_dpath_pmp_4_cfg_w),
    .io_dpath_pmp_4_cfg_r(ptw_io_dpath_pmp_4_cfg_r),
    .io_dpath_pmp_4_addr(ptw_io_dpath_pmp_4_addr),
    .io_dpath_pmp_4_mask(ptw_io_dpath_pmp_4_mask),
    .io_dpath_pmp_5_cfg_l(ptw_io_dpath_pmp_5_cfg_l),
    .io_dpath_pmp_5_cfg_a(ptw_io_dpath_pmp_5_cfg_a),
    .io_dpath_pmp_5_cfg_x(ptw_io_dpath_pmp_5_cfg_x),
    .io_dpath_pmp_5_cfg_w(ptw_io_dpath_pmp_5_cfg_w),
    .io_dpath_pmp_5_cfg_r(ptw_io_dpath_pmp_5_cfg_r),
    .io_dpath_pmp_5_addr(ptw_io_dpath_pmp_5_addr),
    .io_dpath_pmp_5_mask(ptw_io_dpath_pmp_5_mask),
    .io_dpath_pmp_6_cfg_l(ptw_io_dpath_pmp_6_cfg_l),
    .io_dpath_pmp_6_cfg_a(ptw_io_dpath_pmp_6_cfg_a),
    .io_dpath_pmp_6_cfg_x(ptw_io_dpath_pmp_6_cfg_x),
    .io_dpath_pmp_6_cfg_w(ptw_io_dpath_pmp_6_cfg_w),
    .io_dpath_pmp_6_cfg_r(ptw_io_dpath_pmp_6_cfg_r),
    .io_dpath_pmp_6_addr(ptw_io_dpath_pmp_6_addr),
    .io_dpath_pmp_6_mask(ptw_io_dpath_pmp_6_mask),
    .io_dpath_pmp_7_cfg_l(ptw_io_dpath_pmp_7_cfg_l),
    .io_dpath_pmp_7_cfg_a(ptw_io_dpath_pmp_7_cfg_a),
    .io_dpath_pmp_7_cfg_x(ptw_io_dpath_pmp_7_cfg_x),
    .io_dpath_pmp_7_cfg_w(ptw_io_dpath_pmp_7_cfg_w),
    .io_dpath_pmp_7_cfg_r(ptw_io_dpath_pmp_7_cfg_r),
    .io_dpath_pmp_7_addr(ptw_io_dpath_pmp_7_addr),
    .io_dpath_pmp_7_mask(ptw_io_dpath_pmp_7_mask)
  );
  Rocket core (
    .clock(core_clock),
    .reset(core_reset),
    .io_hartid(core_io_hartid),
    .io_interrupts_debug(core_io_interrupts_debug),
    .io_interrupts_mtip(core_io_interrupts_mtip),
    .io_interrupts_msip(core_io_interrupts_msip),
    .io_interrupts_meip(core_io_interrupts_meip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_sfence_valid(core_io_imem_sfence_valid),
    .io_imem_sfence_bits_rs1(core_io_imem_sfence_bits_rs1),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_btb_valid(core_io_imem_resp_bits_btb_valid),
    .io_imem_resp_bits_btb_bits_taken(core_io_imem_resp_bits_btb_bits_taken),
    .io_imem_resp_bits_btb_bits_bridx(core_io_imem_resp_bits_btb_bits_bridx),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_imem_resp_bits_xcpt_pf_inst(core_io_imem_resp_bits_xcpt_pf_inst),
    .io_imem_resp_bits_xcpt_ae_inst(core_io_imem_resp_bits_xcpt_ae_inst),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data_data(core_io_dmem_s1_data_data),
    .io_dmem_s1_data_mask(core_io_dmem_s1_data_mask),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_s2_xcpt_ma_ld(core_io_dmem_s2_xcpt_ma_ld),
    .io_dmem_s2_xcpt_ma_st(core_io_dmem_s2_xcpt_ma_st),
    .io_dmem_s2_xcpt_pf_ld(core_io_dmem_s2_xcpt_pf_ld),
    .io_dmem_s2_xcpt_pf_st(core_io_dmem_s2_xcpt_pf_st),
    .io_dmem_s2_xcpt_ae_ld(core_io_dmem_s2_xcpt_ae_ld),
    .io_dmem_s2_xcpt_ae_st(core_io_dmem_s2_xcpt_ae_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_sfence_valid(core_io_ptw_sfence_valid),
    .io_ptw_sfence_bits_rs1(core_io_ptw_sfence_bits_rs1),
    .io_ptw_status_dprv(core_io_ptw_status_dprv),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_sum(core_io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l(core_io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a(core_io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x(core_io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w(core_io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r(core_io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr(core_io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask(core_io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l(core_io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a(core_io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x(core_io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w(core_io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r(core_io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr(core_io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask(core_io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l(core_io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a(core_io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x(core_io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w(core_io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r(core_io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr(core_io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask(core_io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l(core_io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a(core_io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x(core_io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w(core_io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r(core_io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr(core_io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask(core_io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l(core_io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a(core_io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x(core_io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w(core_io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r(core_io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr(core_io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask(core_io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l(core_io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a(core_io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x(core_io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w(core_io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r(core_io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr(core_io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask(core_io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l(core_io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a(core_io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x(core_io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w(core_io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r(core_io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr(core_io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask(core_io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l(core_io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a(core_io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x(core_io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w(core_io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r(core_io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr(core_io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask(core_io_ptw_pmp_7_mask),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_interrupt(core_io_rocc_interrupt)
  );
  assign io_master_0_a_valid = tileBus_io_out_0_a_valid;
  assign io_master_0_a_bits_opcode = tileBus_io_out_0_a_bits_opcode;
  assign io_master_0_a_bits_param = tileBus_io_out_0_a_bits_param;
  assign io_master_0_a_bits_size = tileBus_io_out_0_a_bits_size;
  assign io_master_0_a_bits_source = tileBus_io_out_0_a_bits_source;
  assign io_master_0_a_bits_address = tileBus_io_out_0_a_bits_address;
  assign io_master_0_a_bits_mask = tileBus_io_out_0_a_bits_mask;
  assign io_master_0_a_bits_data = tileBus_io_out_0_a_bits_data;
  assign io_master_0_d_ready = tileBus_io_out_0_d_ready;
  assign io_slave_0_a_ready = TLFragmenter_io_in_0_a_ready;
  assign io_slave_0_d_valid = TLFragmenter_io_in_0_d_valid;
  assign io_slave_0_d_bits_opcode = TLFragmenter_io_in_0_d_bits_opcode;
  assign io_slave_0_d_bits_param = TLFragmenter_io_in_0_d_bits_param;
  assign io_slave_0_d_bits_size = TLFragmenter_io_in_0_d_bits_size;
  assign io_slave_0_d_bits_source = TLFragmenter_io_in_0_d_bits_source;
  assign io_slave_0_d_bits_sink = TLFragmenter_io_in_0_d_bits_sink;
  assign io_slave_0_d_bits_data = TLFragmenter_io_in_0_d_bits_data;
  assign io_slave_0_d_bits_error = TLFragmenter_io_in_0_d_bits_error;
  assign tileBus_clock = clock;
  assign tileBus_reset = reset;
  assign tileBus_io_in_1_a_valid = frontend_io_tl_out_0_a_valid;
  assign tileBus_io_in_1_a_bits_opcode = frontend_io_tl_out_0_a_bits_opcode;
  assign tileBus_io_in_1_a_bits_param = frontend_io_tl_out_0_a_bits_param;
  assign tileBus_io_in_1_a_bits_size = frontend_io_tl_out_0_a_bits_size;
  assign tileBus_io_in_1_a_bits_source = frontend_io_tl_out_0_a_bits_source;
  assign tileBus_io_in_1_a_bits_address = frontend_io_tl_out_0_a_bits_address;
  assign tileBus_io_in_1_a_bits_mask = frontend_io_tl_out_0_a_bits_mask;
  assign tileBus_io_in_1_a_bits_data = frontend_io_tl_out_0_a_bits_data;
  assign tileBus_io_in_1_d_ready = frontend_io_tl_out_0_d_ready;
  assign tileBus_io_in_0_a_valid = dcache_io_mem_0_a_valid;
  assign tileBus_io_in_0_a_bits_opcode = dcache_io_mem_0_a_bits_opcode;
  assign tileBus_io_in_0_a_bits_param = dcache_io_mem_0_a_bits_param;
  assign tileBus_io_in_0_a_bits_size = dcache_io_mem_0_a_bits_size;
  assign tileBus_io_in_0_a_bits_address = dcache_io_mem_0_a_bits_address;
  assign tileBus_io_in_0_a_bits_mask = dcache_io_mem_0_a_bits_mask;
  assign tileBus_io_in_0_a_bits_data = dcache_io_mem_0_a_bits_data;
  assign tileBus_io_in_0_d_ready = dcache_io_mem_0_d_ready;
  assign tileBus_io_out_0_a_ready = io_master_0_a_ready;
  assign tileBus_io_out_0_d_valid = io_master_0_d_valid;
  assign tileBus_io_out_0_d_bits_opcode = io_master_0_d_bits_opcode;
  assign tileBus_io_out_0_d_bits_size = io_master_0_d_bits_size;
  assign tileBus_io_out_0_d_bits_source = io_master_0_d_bits_source;
  assign tileBus_io_out_0_d_bits_data = io_master_0_d_bits_data;
  assign tileBus_io_out_0_d_bits_error = io_master_0_d_bits_error;
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_cpu_req_valid = dcacheArb_io_mem_req_valid;
  assign dcache_io_cpu_req_bits_addr = dcacheArb_io_mem_req_bits_addr;
  assign dcache_io_cpu_req_bits_tag = dcacheArb_io_mem_req_bits_tag;
  assign dcache_io_cpu_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd;
  assign dcache_io_cpu_req_bits_typ = dcacheArb_io_mem_req_bits_typ;
  assign dcache_io_cpu_req_bits_phys = dcacheArb_io_mem_req_bits_phys;
  assign dcache_io_cpu_s1_kill = dcacheArb_io_mem_s1_kill;
  assign dcache_io_cpu_s1_data_data = dcacheArb_io_mem_s1_data_data;
  assign dcache_io_cpu_s1_data_mask = dcacheArb_io_mem_s1_data_mask;
  assign dcache_io_cpu_invalidate_lr = dcacheArb_io_mem_invalidate_lr;
  assign dcache_io_ptw_resp_valid = ptw_io_requestor_0_resp_valid;
  assign dcache_io_ptw_status_dprv = ptw_io_requestor_0_status_dprv;
  assign dcache_io_ptw_status_prv = ptw_io_requestor_0_status_prv;
  assign dcache_io_ptw_status_mxr = ptw_io_requestor_0_status_mxr;
  assign dcache_io_ptw_status_sum = ptw_io_requestor_0_status_sum;
  assign dcache_io_ptw_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l;
  assign dcache_io_ptw_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a;
  assign dcache_io_ptw_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x;
  assign dcache_io_ptw_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w;
  assign dcache_io_ptw_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r;
  assign dcache_io_ptw_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr;
  assign dcache_io_ptw_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask;
  assign dcache_io_ptw_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l;
  assign dcache_io_ptw_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a;
  assign dcache_io_ptw_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x;
  assign dcache_io_ptw_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w;
  assign dcache_io_ptw_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r;
  assign dcache_io_ptw_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr;
  assign dcache_io_ptw_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask;
  assign dcache_io_ptw_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l;
  assign dcache_io_ptw_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a;
  assign dcache_io_ptw_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x;
  assign dcache_io_ptw_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w;
  assign dcache_io_ptw_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r;
  assign dcache_io_ptw_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr;
  assign dcache_io_ptw_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask;
  assign dcache_io_ptw_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l;
  assign dcache_io_ptw_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a;
  assign dcache_io_ptw_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x;
  assign dcache_io_ptw_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w;
  assign dcache_io_ptw_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r;
  assign dcache_io_ptw_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr;
  assign dcache_io_ptw_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask;
  assign dcache_io_ptw_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l;
  assign dcache_io_ptw_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a;
  assign dcache_io_ptw_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x;
  assign dcache_io_ptw_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w;
  assign dcache_io_ptw_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r;
  assign dcache_io_ptw_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr;
  assign dcache_io_ptw_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask;
  assign dcache_io_ptw_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l;
  assign dcache_io_ptw_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a;
  assign dcache_io_ptw_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x;
  assign dcache_io_ptw_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w;
  assign dcache_io_ptw_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r;
  assign dcache_io_ptw_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr;
  assign dcache_io_ptw_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask;
  assign dcache_io_ptw_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l;
  assign dcache_io_ptw_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a;
  assign dcache_io_ptw_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x;
  assign dcache_io_ptw_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w;
  assign dcache_io_ptw_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r;
  assign dcache_io_ptw_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr;
  assign dcache_io_ptw_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask;
  assign dcache_io_ptw_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l;
  assign dcache_io_ptw_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a;
  assign dcache_io_ptw_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x;
  assign dcache_io_ptw_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w;
  assign dcache_io_ptw_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r;
  assign dcache_io_ptw_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr;
  assign dcache_io_ptw_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask;
  assign dcache_io_mem_0_a_ready = tileBus_io_in_0_a_ready;
  assign dcache_io_mem_0_b_valid = tileBus_io_in_0_b_valid;
  assign dcache_io_mem_0_b_bits_param = tileBus_io_in_0_b_bits_param;
  assign dcache_io_mem_0_b_bits_address = tileBus_io_in_0_b_bits_address;
  assign dcache_io_mem_0_c_ready = tileBus_io_in_0_c_ready;
  assign dcache_io_mem_0_d_valid = tileBus_io_in_0_d_valid;
  assign dcache_io_mem_0_d_bits_opcode = tileBus_io_in_0_d_bits_opcode;
  assign dcache_io_mem_0_d_bits_size = tileBus_io_in_0_d_bits_size;
  assign dcache_io_mem_0_d_bits_source = tileBus_io_in_0_d_bits_source;
  assign dcache_io_mem_0_d_bits_data = tileBus_io_in_0_d_bits_data;
  assign dcache_io_mem_0_e_ready = tileBus_io_in_0_e_ready;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_tl_out_0_a_ready = tileBus_io_in_1_a_ready;
  assign frontend_io_tl_out_0_d_valid = tileBus_io_in_1_d_valid;
  assign frontend_io_tl_out_0_d_bits_opcode = tileBus_io_in_1_d_bits_opcode;
  assign frontend_io_tl_out_0_d_bits_size = tileBus_io_in_1_d_bits_size;
  assign frontend_io_tl_out_0_d_bits_data = tileBus_io_in_1_d_bits_data;
  assign frontend_io_tl_out_0_d_bits_error = tileBus_io_in_1_d_bits_error;
  assign frontend_io_cpu_req_valid = core_io_imem_req_valid;
  assign frontend_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign frontend_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
  assign frontend_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign frontend_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign frontend_io_ptw_resp_valid = ptw_io_requestor_1_resp_valid;
  assign frontend_io_ptw_status_dprv = ptw_io_requestor_1_status_dprv;
  assign frontend_io_ptw_status_prv = ptw_io_requestor_1_status_prv;
  assign frontend_io_ptw_status_mxr = ptw_io_requestor_1_status_mxr;
  assign frontend_io_ptw_status_sum = ptw_io_requestor_1_status_sum;
  assign frontend_io_ptw_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l;
  assign frontend_io_ptw_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a;
  assign frontend_io_ptw_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x;
  assign frontend_io_ptw_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w;
  assign frontend_io_ptw_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r;
  assign frontend_io_ptw_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr;
  assign frontend_io_ptw_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask;
  assign frontend_io_ptw_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l;
  assign frontend_io_ptw_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a;
  assign frontend_io_ptw_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x;
  assign frontend_io_ptw_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w;
  assign frontend_io_ptw_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r;
  assign frontend_io_ptw_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr;
  assign frontend_io_ptw_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask;
  assign frontend_io_ptw_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l;
  assign frontend_io_ptw_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a;
  assign frontend_io_ptw_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x;
  assign frontend_io_ptw_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w;
  assign frontend_io_ptw_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r;
  assign frontend_io_ptw_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr;
  assign frontend_io_ptw_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask;
  assign frontend_io_ptw_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l;
  assign frontend_io_ptw_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a;
  assign frontend_io_ptw_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x;
  assign frontend_io_ptw_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w;
  assign frontend_io_ptw_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r;
  assign frontend_io_ptw_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr;
  assign frontend_io_ptw_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask;
  assign frontend_io_ptw_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l;
  assign frontend_io_ptw_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a;
  assign frontend_io_ptw_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x;
  assign frontend_io_ptw_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w;
  assign frontend_io_ptw_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r;
  assign frontend_io_ptw_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr;
  assign frontend_io_ptw_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask;
  assign frontend_io_ptw_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l;
  assign frontend_io_ptw_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a;
  assign frontend_io_ptw_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x;
  assign frontend_io_ptw_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w;
  assign frontend_io_ptw_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r;
  assign frontend_io_ptw_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr;
  assign frontend_io_ptw_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask;
  assign frontend_io_ptw_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l;
  assign frontend_io_ptw_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a;
  assign frontend_io_ptw_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x;
  assign frontend_io_ptw_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w;
  assign frontend_io_ptw_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r;
  assign frontend_io_ptw_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr;
  assign frontend_io_ptw_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask;
  assign frontend_io_ptw_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l;
  assign frontend_io_ptw_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a;
  assign frontend_io_ptw_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x;
  assign frontend_io_ptw_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w;
  assign frontend_io_ptw_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r;
  assign frontend_io_ptw_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr;
  assign frontend_io_ptw_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask;
  assign frontend_io_resetVector = io_resetVector;
  assign ScratchpadSlavePort_clock = clock;
  assign ScratchpadSlavePort_reset = reset;
  assign ScratchpadSlavePort_io_tl_in_0_a_valid = TLFragmenter_io_out_0_a_valid;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_opcode = TLFragmenter_io_out_0_a_bits_opcode;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_param = TLFragmenter_io_out_0_a_bits_param;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_size = TLFragmenter_io_out_0_a_bits_size;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_source = TLFragmenter_io_out_0_a_bits_source;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_address = TLFragmenter_io_out_0_a_bits_address;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_mask = TLFragmenter_io_out_0_a_bits_mask;
  assign ScratchpadSlavePort_io_tl_in_0_a_bits_data = TLFragmenter_io_out_0_a_bits_data;
  assign ScratchpadSlavePort_io_tl_in_0_d_ready = TLFragmenter_io_out_0_d_ready;
  assign ScratchpadSlavePort_io_dmem_req_ready = dcacheArb_io_requestor_0_req_ready;
  assign ScratchpadSlavePort_io_dmem_s2_nack = dcacheArb_io_requestor_0_s2_nack;
  assign ScratchpadSlavePort_io_dmem_resp_valid = dcacheArb_io_requestor_0_resp_valid;
  assign ScratchpadSlavePort_io_dmem_resp_bits_data_raw = dcacheArb_io_requestor_0_resp_bits_data_raw;
  assign TLFragmenter_clock = clock;
  assign TLFragmenter_reset = reset;
  assign TLFragmenter_io_in_0_a_valid = io_slave_0_a_valid;
  assign TLFragmenter_io_in_0_a_bits_opcode = io_slave_0_a_bits_opcode;
  assign TLFragmenter_io_in_0_a_bits_param = io_slave_0_a_bits_param;
  assign TLFragmenter_io_in_0_a_bits_size = io_slave_0_a_bits_size;
  assign TLFragmenter_io_in_0_a_bits_source = io_slave_0_a_bits_source;
  assign TLFragmenter_io_in_0_a_bits_address = io_slave_0_a_bits_address;
  assign TLFragmenter_io_in_0_a_bits_mask = io_slave_0_a_bits_mask;
  assign TLFragmenter_io_in_0_a_bits_data = io_slave_0_a_bits_data;
  assign TLFragmenter_io_in_0_d_ready = io_slave_0_d_ready;
  assign TLFragmenter_io_out_0_a_ready = ScratchpadSlavePort_io_tl_in_0_a_ready;
  assign TLFragmenter_io_out_0_d_valid = ScratchpadSlavePort_io_tl_in_0_d_valid;
  assign TLFragmenter_io_out_0_d_bits_opcode = ScratchpadSlavePort_io_tl_in_0_d_bits_opcode;
  assign TLFragmenter_io_out_0_d_bits_param = ScratchpadSlavePort_io_tl_in_0_d_bits_param;
  assign TLFragmenter_io_out_0_d_bits_size = ScratchpadSlavePort_io_tl_in_0_d_bits_size;
  assign TLFragmenter_io_out_0_d_bits_source = ScratchpadSlavePort_io_tl_in_0_d_bits_source;
  assign TLFragmenter_io_out_0_d_bits_sink = ScratchpadSlavePort_io_tl_in_0_d_bits_sink;
  assign TLFragmenter_io_out_0_d_bits_data = ScratchpadSlavePort_io_tl_in_0_d_bits_data;
  assign TLFragmenter_io_out_0_d_bits_error = ScratchpadSlavePort_io_tl_in_0_d_bits_error;
  assign dcacheArb_clock = clock;
  assign dcacheArb_io_requestor_0_req_valid = ScratchpadSlavePort_io_dmem_req_valid;
  assign dcacheArb_io_requestor_0_req_bits_addr = ScratchpadSlavePort_io_dmem_req_bits_addr;
  assign dcacheArb_io_requestor_0_req_bits_tag = ScratchpadSlavePort_io_dmem_req_bits_tag;
  assign dcacheArb_io_requestor_0_req_bits_cmd = ScratchpadSlavePort_io_dmem_req_bits_cmd;
  assign dcacheArb_io_requestor_0_req_bits_typ = ScratchpadSlavePort_io_dmem_req_bits_typ;
  assign dcacheArb_io_requestor_0_req_bits_phys = ScratchpadSlavePort_io_dmem_req_bits_phys;
  assign dcacheArb_io_requestor_0_s1_kill = ScratchpadSlavePort_io_dmem_s1_kill;
  assign dcacheArb_io_requestor_0_s1_data_data = ScratchpadSlavePort_io_dmem_s1_data_data;
  assign dcacheArb_io_requestor_0_s1_data_mask = ScratchpadSlavePort_io_dmem_s1_data_mask;
  assign dcacheArb_io_requestor_0_invalidate_lr = ScratchpadSlavePort_io_dmem_invalidate_lr;
  assign dcacheArb_io_requestor_1_req_valid = core_io_dmem_req_valid;
  assign dcacheArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcacheArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcacheArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcacheArb_io_requestor_1_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcacheArb_io_requestor_1_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcacheArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill;
  assign dcacheArb_io_requestor_1_s1_data_data = core_io_dmem_s1_data_data;
  assign dcacheArb_io_requestor_1_s1_data_mask = core_io_dmem_s1_data_mask;
  assign dcacheArb_io_requestor_1_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcacheArb_io_mem_req_ready = dcache_io_cpu_req_ready;
  assign dcacheArb_io_mem_s2_nack = dcache_io_cpu_s2_nack;
  assign dcacheArb_io_mem_resp_valid = dcache_io_cpu_resp_valid;
  assign dcacheArb_io_mem_resp_bits_tag = dcache_io_cpu_resp_bits_tag;
  assign dcacheArb_io_mem_resp_bits_data = dcache_io_cpu_resp_bits_data;
  assign dcacheArb_io_mem_resp_bits_replay = dcache_io_cpu_resp_bits_replay;
  assign dcacheArb_io_mem_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data;
  assign dcacheArb_io_mem_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass;
  assign dcacheArb_io_mem_resp_bits_data_raw = dcache_io_cpu_resp_bits_data_raw;
  assign dcacheArb_io_mem_replay_next = dcache_io_cpu_replay_next;
  assign dcacheArb_io_mem_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld;
  assign dcacheArb_io_mem_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st;
  assign dcacheArb_io_mem_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld;
  assign dcacheArb_io_mem_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st;
  assign dcacheArb_io_mem_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld;
  assign dcacheArb_io_mem_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st;
  assign dcacheArb_io_mem_ordered = dcache_io_cpu_ordered;
  assign ptw_clock = clock;
  assign ptw_reset = reset;
  assign ptw_io_requestor_0_req_valid = dcache_io_ptw_req_valid;
  assign ptw_io_requestor_0_req_bits_addr = dcache_io_ptw_req_bits_addr;
  assign ptw_io_requestor_1_req_valid = frontend_io_ptw_req_valid;
  assign ptw_io_requestor_1_req_bits_addr = frontend_io_ptw_req_bits_addr;
  assign ptw_io_mem_req_ready = 1'h0;
  assign ptw_io_mem_s2_nack = 1'h0;
  assign ptw_io_mem_resp_valid = 1'h0;
  assign ptw_io_mem_resp_bits_data = 32'h0;
  assign ptw_io_mem_s2_xcpt_ae_ld = 1'h0;
  assign ptw_io_dpath_ptbr_ppn = core_io_ptw_ptbr_ppn;
  assign ptw_io_dpath_sfence_valid = core_io_ptw_sfence_valid;
  assign ptw_io_dpath_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1;
  assign ptw_io_dpath_status_dprv = core_io_ptw_status_dprv;
  assign ptw_io_dpath_status_prv = core_io_ptw_status_prv;
  assign ptw_io_dpath_status_mxr = core_io_ptw_status_mxr;
  assign ptw_io_dpath_status_sum = core_io_ptw_status_sum;
  assign ptw_io_dpath_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l;
  assign ptw_io_dpath_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a;
  assign ptw_io_dpath_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x;
  assign ptw_io_dpath_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w;
  assign ptw_io_dpath_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r;
  assign ptw_io_dpath_pmp_0_addr = core_io_ptw_pmp_0_addr;
  assign ptw_io_dpath_pmp_0_mask = core_io_ptw_pmp_0_mask;
  assign ptw_io_dpath_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l;
  assign ptw_io_dpath_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a;
  assign ptw_io_dpath_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x;
  assign ptw_io_dpath_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w;
  assign ptw_io_dpath_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r;
  assign ptw_io_dpath_pmp_1_addr = core_io_ptw_pmp_1_addr;
  assign ptw_io_dpath_pmp_1_mask = core_io_ptw_pmp_1_mask;
  assign ptw_io_dpath_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l;
  assign ptw_io_dpath_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a;
  assign ptw_io_dpath_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x;
  assign ptw_io_dpath_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w;
  assign ptw_io_dpath_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r;
  assign ptw_io_dpath_pmp_2_addr = core_io_ptw_pmp_2_addr;
  assign ptw_io_dpath_pmp_2_mask = core_io_ptw_pmp_2_mask;
  assign ptw_io_dpath_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l;
  assign ptw_io_dpath_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a;
  assign ptw_io_dpath_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x;
  assign ptw_io_dpath_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w;
  assign ptw_io_dpath_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r;
  assign ptw_io_dpath_pmp_3_addr = core_io_ptw_pmp_3_addr;
  assign ptw_io_dpath_pmp_3_mask = core_io_ptw_pmp_3_mask;
  assign ptw_io_dpath_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l;
  assign ptw_io_dpath_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a;
  assign ptw_io_dpath_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x;
  assign ptw_io_dpath_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w;
  assign ptw_io_dpath_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r;
  assign ptw_io_dpath_pmp_4_addr = core_io_ptw_pmp_4_addr;
  assign ptw_io_dpath_pmp_4_mask = core_io_ptw_pmp_4_mask;
  assign ptw_io_dpath_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l;
  assign ptw_io_dpath_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a;
  assign ptw_io_dpath_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x;
  assign ptw_io_dpath_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w;
  assign ptw_io_dpath_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r;
  assign ptw_io_dpath_pmp_5_addr = core_io_ptw_pmp_5_addr;
  assign ptw_io_dpath_pmp_5_mask = core_io_ptw_pmp_5_mask;
  assign ptw_io_dpath_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l;
  assign ptw_io_dpath_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a;
  assign ptw_io_dpath_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x;
  assign ptw_io_dpath_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w;
  assign ptw_io_dpath_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r;
  assign ptw_io_dpath_pmp_6_addr = core_io_ptw_pmp_6_addr;
  assign ptw_io_dpath_pmp_6_mask = core_io_ptw_pmp_6_mask;
  assign ptw_io_dpath_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l;
  assign ptw_io_dpath_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a;
  assign ptw_io_dpath_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x;
  assign ptw_io_dpath_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w;
  assign ptw_io_dpath_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r;
  assign ptw_io_dpath_pmp_7_addr = core_io_ptw_pmp_7_addr;
  assign ptw_io_dpath_pmp_7_mask = core_io_ptw_pmp_7_mask;
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_hartid = io_hartid;
  assign core_io_interrupts_debug = io_interrupts_0_0;
  assign core_io_interrupts_mtip = io_interrupts_0_2;
  assign core_io_interrupts_msip = io_interrupts_0_1;
  assign core_io_interrupts_meip = io_interrupts_0_3;
  assign core_io_imem_resp_valid = frontend_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_btb_valid = frontend_io_cpu_resp_bits_btb_valid;
  assign core_io_imem_resp_bits_btb_bits_taken = frontend_io_cpu_resp_bits_btb_bits_taken;
  assign core_io_imem_resp_bits_btb_bits_bridx = frontend_io_cpu_resp_bits_btb_bits_bridx;
  assign core_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data = frontend_io_cpu_resp_bits_data;
  assign core_io_imem_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst;
  assign core_io_imem_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst;
  assign core_io_imem_resp_bits_replay = frontend_io_cpu_resp_bits_replay;
  assign core_io_dmem_req_ready = dcacheArb_io_requestor_1_req_ready;
  assign core_io_dmem_s2_nack = dcacheArb_io_requestor_1_s2_nack;
  assign core_io_dmem_resp_valid = dcacheArb_io_requestor_1_resp_valid;
  assign core_io_dmem_resp_bits_tag = dcacheArb_io_requestor_1_resp_bits_tag;
  assign core_io_dmem_resp_bits_data = dcacheArb_io_requestor_1_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcacheArb_io_requestor_1_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcacheArb_io_requestor_1_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcacheArb_io_requestor_1_resp_bits_data_word_bypass;
  assign core_io_dmem_replay_next = dcacheArb_io_requestor_1_replay_next;
  assign core_io_dmem_s2_xcpt_ma_ld = dcacheArb_io_requestor_1_s2_xcpt_ma_ld;
  assign core_io_dmem_s2_xcpt_ma_st = dcacheArb_io_requestor_1_s2_xcpt_ma_st;
  assign core_io_dmem_s2_xcpt_pf_ld = dcacheArb_io_requestor_1_s2_xcpt_pf_ld;
  assign core_io_dmem_s2_xcpt_pf_st = dcacheArb_io_requestor_1_s2_xcpt_pf_st;
  assign core_io_dmem_s2_xcpt_ae_ld = dcacheArb_io_requestor_1_s2_xcpt_ae_ld;
  assign core_io_dmem_s2_xcpt_ae_st = dcacheArb_io_requestor_1_s2_xcpt_ae_st;
  assign core_io_dmem_ordered = dcacheArb_io_requestor_1_ordered;
  assign core_io_fpu_store_data = 32'h0;
  assign core_io_fpu_toint_data = 32'h0;
  assign core_io_fpu_nack_mem = 1'h0;
  assign core_io_fpu_dec_wen = 1'h0;
  assign core_io_fpu_dec_ren1 = 1'h0;
  assign core_io_fpu_dec_ren2 = 1'h0;
  assign core_io_fpu_dec_ren3 = 1'h0;
  assign core_io_rocc_cmd_ready = 1'h0;
  assign core_io_rocc_interrupt = 1'h0;
endmodule
module IntXbar_intXbar(
  input   io_in_1_0,
  input   io_in_1_1,
  input   io_in_1_2,
  input   io_in_0_0,
  output  io_out_0_0,
  output  io_out_0_1,
  output  io_out_0_2,
  output  io_out_0_3
);
  assign io_out_0_0 = io_in_0_0;
  assign io_out_0_1 = io_in_1_0;
  assign io_out_0_2 = io_in_1_1;
  assign io_out_0_3 = io_in_1_2;
endmodule
module IntXing_xing(
  input   clock,
  input   io_in_0_0,
  output  io_out_0_0
);
  reg  _T_19_0;
  reg [31:0] _RAND_0;
  reg  _T_37_0;
  reg [31:0] _RAND_1;
  reg  _T_63_0;
  reg [31:0] _RAND_2;
  reg  _T_97_0;
  reg [31:0] _RAND_3;
  assign io_out_0_0 = _T_97_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_19_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_37_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_63_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_97_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_19_0 <= io_in_0_0;
    _T_37_0 <= _T_19_0;
    _T_63_0 <= _T_37_0;
    _T_97_0 <= _T_63_0;
  end
endmodule
module SyncRocketTile_tile(
  input         clock,
  input         reset,
  input         io_master_0_a_ready,
  output        io_master_0_a_valid,
  output [2:0]  io_master_0_a_bits_opcode,
  output [2:0]  io_master_0_a_bits_param,
  output [3:0]  io_master_0_a_bits_size,
  output        io_master_0_a_bits_source,
  output [31:0] io_master_0_a_bits_address,
  output [3:0]  io_master_0_a_bits_mask,
  output [31:0] io_master_0_a_bits_data,
  output        io_master_0_d_ready,
  input         io_master_0_d_valid,
  input  [2:0]  io_master_0_d_bits_opcode,
  input  [3:0]  io_master_0_d_bits_size,
  input         io_master_0_d_bits_source,
  input  [31:0] io_master_0_d_bits_data,
  input         io_master_0_d_bits_error,
  output        io_slave_0_a_ready,
  input         io_slave_0_a_valid,
  input  [2:0]  io_slave_0_a_bits_opcode,
  input  [2:0]  io_slave_0_a_bits_param,
  input  [2:0]  io_slave_0_a_bits_size,
  input  [4:0]  io_slave_0_a_bits_source,
  input  [31:0] io_slave_0_a_bits_address,
  input  [3:0]  io_slave_0_a_bits_mask,
  input  [31:0] io_slave_0_a_bits_data,
  input         io_slave_0_d_ready,
  output        io_slave_0_d_valid,
  output [2:0]  io_slave_0_d_bits_opcode,
  output [1:0]  io_slave_0_d_bits_param,
  output [2:0]  io_slave_0_d_bits_size,
  output [4:0]  io_slave_0_d_bits_source,
  output        io_slave_0_d_bits_sink,
  output [31:0] io_slave_0_d_bits_data,
  output        io_slave_0_d_bits_error,
  input         io_asyncInterrupts_0_0,
  input         io_periphInterrupts_0_0,
  input         io_periphInterrupts_0_1,
  input         io_periphInterrupts_0_2,
  input         io_hartid,
  input  [31:0] io_resetVector
);
  wire  rocket_clock;
  wire  rocket_reset;
  wire  rocket_io_master_0_a_ready;
  wire  rocket_io_master_0_a_valid;
  wire [2:0] rocket_io_master_0_a_bits_opcode;
  wire [2:0] rocket_io_master_0_a_bits_param;
  wire [3:0] rocket_io_master_0_a_bits_size;
  wire  rocket_io_master_0_a_bits_source;
  wire [31:0] rocket_io_master_0_a_bits_address;
  wire [3:0] rocket_io_master_0_a_bits_mask;
  wire [31:0] rocket_io_master_0_a_bits_data;
  wire  rocket_io_master_0_d_ready;
  wire  rocket_io_master_0_d_valid;
  wire [2:0] rocket_io_master_0_d_bits_opcode;
  wire [3:0] rocket_io_master_0_d_bits_size;
  wire  rocket_io_master_0_d_bits_source;
  wire [31:0] rocket_io_master_0_d_bits_data;
  wire  rocket_io_master_0_d_bits_error;
  wire  rocket_io_slave_0_a_ready;
  wire  rocket_io_slave_0_a_valid;
  wire [2:0] rocket_io_slave_0_a_bits_opcode;
  wire [2:0] rocket_io_slave_0_a_bits_param;
  wire [2:0] rocket_io_slave_0_a_bits_size;
  wire [4:0] rocket_io_slave_0_a_bits_source;
  wire [31:0] rocket_io_slave_0_a_bits_address;
  wire [3:0] rocket_io_slave_0_a_bits_mask;
  wire [31:0] rocket_io_slave_0_a_bits_data;
  wire  rocket_io_slave_0_d_ready;
  wire  rocket_io_slave_0_d_valid;
  wire [2:0] rocket_io_slave_0_d_bits_opcode;
  wire [1:0] rocket_io_slave_0_d_bits_param;
  wire [2:0] rocket_io_slave_0_d_bits_size;
  wire [4:0] rocket_io_slave_0_d_bits_source;
  wire  rocket_io_slave_0_d_bits_sink;
  wire [31:0] rocket_io_slave_0_d_bits_data;
  wire  rocket_io_slave_0_d_bits_error;
  wire  rocket_io_hartid;
  wire [31:0] rocket_io_resetVector;
  wire  rocket_io_interrupts_0_0;
  wire  rocket_io_interrupts_0_1;
  wire  rocket_io_interrupts_0_2;
  wire  rocket_io_interrupts_0_3;
  wire  intXbar_io_in_1_0;
  wire  intXbar_io_in_1_1;
  wire  intXbar_io_in_1_2;
  wire  intXbar_io_in_0_0;
  wire  intXbar_io_out_0_0;
  wire  intXbar_io_out_0_1;
  wire  intXbar_io_out_0_2;
  wire  intXbar_io_out_0_3;
  wire  xing_clock;
  wire  xing_io_in_0_0;
  wire  xing_io_out_0_0;
  RocketTile_rocket rocket (
    .clock(rocket_clock),
    .reset(rocket_reset),
    .io_master_0_a_ready(rocket_io_master_0_a_ready),
    .io_master_0_a_valid(rocket_io_master_0_a_valid),
    .io_master_0_a_bits_opcode(rocket_io_master_0_a_bits_opcode),
    .io_master_0_a_bits_param(rocket_io_master_0_a_bits_param),
    .io_master_0_a_bits_size(rocket_io_master_0_a_bits_size),
    .io_master_0_a_bits_source(rocket_io_master_0_a_bits_source),
    .io_master_0_a_bits_address(rocket_io_master_0_a_bits_address),
    .io_master_0_a_bits_mask(rocket_io_master_0_a_bits_mask),
    .io_master_0_a_bits_data(rocket_io_master_0_a_bits_data),
    .io_master_0_d_ready(rocket_io_master_0_d_ready),
    .io_master_0_d_valid(rocket_io_master_0_d_valid),
    .io_master_0_d_bits_opcode(rocket_io_master_0_d_bits_opcode),
    .io_master_0_d_bits_size(rocket_io_master_0_d_bits_size),
    .io_master_0_d_bits_source(rocket_io_master_0_d_bits_source),
    .io_master_0_d_bits_data(rocket_io_master_0_d_bits_data),
    .io_master_0_d_bits_error(rocket_io_master_0_d_bits_error),
    .io_slave_0_a_ready(rocket_io_slave_0_a_ready),
    .io_slave_0_a_valid(rocket_io_slave_0_a_valid),
    .io_slave_0_a_bits_opcode(rocket_io_slave_0_a_bits_opcode),
    .io_slave_0_a_bits_param(rocket_io_slave_0_a_bits_param),
    .io_slave_0_a_bits_size(rocket_io_slave_0_a_bits_size),
    .io_slave_0_a_bits_source(rocket_io_slave_0_a_bits_source),
    .io_slave_0_a_bits_address(rocket_io_slave_0_a_bits_address),
    .io_slave_0_a_bits_mask(rocket_io_slave_0_a_bits_mask),
    .io_slave_0_a_bits_data(rocket_io_slave_0_a_bits_data),
    .io_slave_0_d_ready(rocket_io_slave_0_d_ready),
    .io_slave_0_d_valid(rocket_io_slave_0_d_valid),
    .io_slave_0_d_bits_opcode(rocket_io_slave_0_d_bits_opcode),
    .io_slave_0_d_bits_param(rocket_io_slave_0_d_bits_param),
    .io_slave_0_d_bits_size(rocket_io_slave_0_d_bits_size),
    .io_slave_0_d_bits_source(rocket_io_slave_0_d_bits_source),
    .io_slave_0_d_bits_sink(rocket_io_slave_0_d_bits_sink),
    .io_slave_0_d_bits_data(rocket_io_slave_0_d_bits_data),
    .io_slave_0_d_bits_error(rocket_io_slave_0_d_bits_error),
    .io_hartid(rocket_io_hartid),
    .io_resetVector(rocket_io_resetVector),
    .io_interrupts_0_0(rocket_io_interrupts_0_0),
    .io_interrupts_0_1(rocket_io_interrupts_0_1),
    .io_interrupts_0_2(rocket_io_interrupts_0_2),
    .io_interrupts_0_3(rocket_io_interrupts_0_3)
  );
  IntXbar_intXbar intXbar (
    .io_in_1_0(intXbar_io_in_1_0),
    .io_in_1_1(intXbar_io_in_1_1),
    .io_in_1_2(intXbar_io_in_1_2),
    .io_in_0_0(intXbar_io_in_0_0),
    .io_out_0_0(intXbar_io_out_0_0),
    .io_out_0_1(intXbar_io_out_0_1),
    .io_out_0_2(intXbar_io_out_0_2),
    .io_out_0_3(intXbar_io_out_0_3)
  );
  IntXing_xing xing (
    .clock(xing_clock),
    .io_in_0_0(xing_io_in_0_0),
    .io_out_0_0(xing_io_out_0_0)
  );
  assign io_master_0_a_valid = rocket_io_master_0_a_valid;
  assign io_master_0_a_bits_opcode = rocket_io_master_0_a_bits_opcode;
  assign io_master_0_a_bits_param = rocket_io_master_0_a_bits_param;
  assign io_master_0_a_bits_size = rocket_io_master_0_a_bits_size;
  assign io_master_0_a_bits_source = rocket_io_master_0_a_bits_source;
  assign io_master_0_a_bits_address = rocket_io_master_0_a_bits_address;
  assign io_master_0_a_bits_mask = rocket_io_master_0_a_bits_mask;
  assign io_master_0_a_bits_data = rocket_io_master_0_a_bits_data;
  assign io_master_0_d_ready = rocket_io_master_0_d_ready;
  assign io_slave_0_a_ready = rocket_io_slave_0_a_ready;
  assign io_slave_0_d_valid = rocket_io_slave_0_d_valid;
  assign io_slave_0_d_bits_opcode = rocket_io_slave_0_d_bits_opcode;
  assign io_slave_0_d_bits_param = rocket_io_slave_0_d_bits_param;
  assign io_slave_0_d_bits_size = rocket_io_slave_0_d_bits_size;
  assign io_slave_0_d_bits_source = rocket_io_slave_0_d_bits_source;
  assign io_slave_0_d_bits_sink = rocket_io_slave_0_d_bits_sink;
  assign io_slave_0_d_bits_data = rocket_io_slave_0_d_bits_data;
  assign io_slave_0_d_bits_error = rocket_io_slave_0_d_bits_error;
  assign rocket_clock = clock;
  assign rocket_reset = reset;
  assign rocket_io_master_0_a_ready = io_master_0_a_ready;
  assign rocket_io_master_0_d_valid = io_master_0_d_valid;
  assign rocket_io_master_0_d_bits_opcode = io_master_0_d_bits_opcode;
  assign rocket_io_master_0_d_bits_size = io_master_0_d_bits_size;
  assign rocket_io_master_0_d_bits_source = io_master_0_d_bits_source;
  assign rocket_io_master_0_d_bits_data = io_master_0_d_bits_data;
  assign rocket_io_master_0_d_bits_error = io_master_0_d_bits_error;
  assign rocket_io_slave_0_a_valid = io_slave_0_a_valid;
  assign rocket_io_slave_0_a_bits_opcode = io_slave_0_a_bits_opcode;
  assign rocket_io_slave_0_a_bits_param = io_slave_0_a_bits_param;
  assign rocket_io_slave_0_a_bits_size = io_slave_0_a_bits_size;
  assign rocket_io_slave_0_a_bits_source = io_slave_0_a_bits_source;
  assign rocket_io_slave_0_a_bits_address = io_slave_0_a_bits_address;
  assign rocket_io_slave_0_a_bits_mask = io_slave_0_a_bits_mask;
  assign rocket_io_slave_0_a_bits_data = io_slave_0_a_bits_data;
  assign rocket_io_slave_0_d_ready = io_slave_0_d_ready;
  assign rocket_io_hartid = io_hartid;
  assign rocket_io_resetVector = io_resetVector;
  assign rocket_io_interrupts_0_0 = intXbar_io_out_0_0;
  assign rocket_io_interrupts_0_1 = intXbar_io_out_0_1;
  assign rocket_io_interrupts_0_2 = intXbar_io_out_0_2;
  assign rocket_io_interrupts_0_3 = intXbar_io_out_0_3;
  assign intXbar_io_in_1_0 = io_periphInterrupts_0_0;
  assign intXbar_io_in_1_1 = io_periphInterrupts_0_1;
  assign intXbar_io_in_1_2 = io_periphInterrupts_0_2;
  assign intXbar_io_in_0_0 = xing_io_out_0_0;
  assign xing_clock = clock;
  assign xing_io_in_0_0 = io_asyncInterrupts_0_0;
endmodule
module Queue_9(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input         io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output        io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_43_data;
  wire  ram_opcode__T_43_addr;
  wire [2:0] ram_opcode__T_29_data;
  wire  ram_opcode__T_29_addr;
  wire  ram_opcode__T_29_mask;
  wire  ram_opcode__T_29_en;
  reg [2:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_43_data;
  wire  ram_param__T_43_addr;
  wire [2:0] ram_param__T_29_data;
  wire  ram_param__T_29_addr;
  wire  ram_param__T_29_mask;
  wire  ram_param__T_29_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [3:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg  ram_source [0:1];
  reg [31:0] _RAND_3;
  wire  ram_source__T_43_data;
  wire  ram_source__T_43_addr;
  wire  ram_source__T_29_data;
  wire  ram_source__T_29_addr;
  wire  ram_source__T_29_mask;
  wire  ram_source__T_29_en;
  reg [31:0] ram_address [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_43_data;
  wire  ram_address__T_43_addr;
  wire [31:0] ram_address__T_29_data;
  wire  ram_address__T_29_addr;
  wire  ram_address__T_29_mask;
  wire  ram_address__T_29_en;
  reg [3:0] ram_mask [0:1];
  reg [31:0] _RAND_5;
  wire [3:0] ram_mask__T_43_data;
  wire  ram_mask__T_43_addr;
  wire [3:0] ram_mask__T_29_data;
  wire  ram_mask__T_29_addr;
  wire  ram_mask__T_29_mask;
  wire  ram_mask__T_29_en;
  reg [31:0] ram_data [0:1];
  reg [31:0] _RAND_6;
  wire [31:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [31:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg  value;
  reg [31:0] _RAND_7;
  reg  value_1;
  reg [31:0] _RAND_8;
  reg  maybe_full;
  reg [31:0] _RAND_9;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_10;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_11;
  wire  _T_38;
  wire  _GEN_12;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_opcode = ram_opcode__T_43_data;
  assign io_deq_bits_param = ram_param__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_source = ram_source__T_43_data;
  assign io_deq_bits_address = ram_address__T_43_data;
  assign io_deq_bits_mask = ram_mask__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign ram_opcode__T_43_addr = value_1;
  assign ram_opcode__T_43_data = ram_opcode[ram_opcode__T_43_addr];
  assign ram_opcode__T_29_data = io_enq_bits_opcode;
  assign ram_opcode__T_29_addr = value;
  assign ram_opcode__T_29_mask = _T_25;
  assign ram_opcode__T_29_en = _T_25;
  assign ram_param__T_43_addr = value_1;
  assign ram_param__T_43_data = ram_param[ram_param__T_43_addr];
  assign ram_param__T_29_data = io_enq_bits_param;
  assign ram_param__T_29_addr = value;
  assign ram_param__T_29_mask = _T_25;
  assign ram_param__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_source__T_43_addr = value_1;
  assign ram_source__T_43_data = ram_source[ram_source__T_43_addr];
  assign ram_source__T_29_data = io_enq_bits_source;
  assign ram_source__T_29_addr = value;
  assign ram_source__T_29_mask = _T_25;
  assign ram_source__T_29_en = _T_25;
  assign ram_address__T_43_addr = value_1;
  assign ram_address__T_43_data = ram_address[ram_address__T_43_addr];
  assign ram_address__T_29_data = io_enq_bits_address;
  assign ram_address__T_29_addr = value;
  assign ram_address__T_29_mask = _T_25;
  assign ram_address__T_29_en = _T_25;
  assign ram_mask__T_43_addr = value_1;
  assign ram_mask__T_43_data = ram_mask[ram_mask__T_43_addr];
  assign ram_mask__T_29_data = io_enq_bits_mask;
  assign ram_mask__T_29_addr = value;
  assign ram_mask__T_29_mask = _T_25;
  assign ram_mask__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_10 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_11 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_12 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_29_en & ram_opcode__T_29_mask) begin
      ram_opcode[ram_opcode__T_29_addr] <= ram_opcode__T_29_data;
    end
    if(ram_param__T_29_en & ram_param__T_29_mask) begin
      ram_param[ram_param__T_29_addr] <= ram_param__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_source__T_29_en & ram_source__T_29_mask) begin
      ram_source[ram_source__T_29_addr] <= ram_source__T_29_data;
    end
    if(ram_address__T_29_en & ram_address__T_29_mask) begin
      ram_address[ram_address__T_29_addr] <= ram_address__T_29_data;
    end
    if(ram_mask__T_29_en & ram_mask__T_29_mask) begin
      ram_mask[ram_mask__T_29_addr] <= ram_mask__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_10(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [3:0]  io_enq_bits_size,
  input         io_enq_bits_source,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [3:0]  io_deq_bits_size,
  output        io_deq_bits_source,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_43_data;
  wire  ram_opcode__T_43_addr;
  wire [2:0] ram_opcode__T_29_data;
  wire  ram_opcode__T_29_addr;
  wire  ram_opcode__T_29_mask;
  wire  ram_opcode__T_29_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [3:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg  ram_source [0:1];
  reg [31:0] _RAND_2;
  wire  ram_source__T_43_data;
  wire  ram_source__T_43_addr;
  wire  ram_source__T_29_data;
  wire  ram_source__T_29_addr;
  wire  ram_source__T_29_mask;
  wire  ram_source__T_29_en;
  reg [31:0] ram_data [0:1];
  reg [31:0] _RAND_3;
  wire [31:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [31:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg  ram_error [0:1];
  reg [31:0] _RAND_4;
  wire  ram_error__T_43_data;
  wire  ram_error__T_43_addr;
  wire  ram_error__T_29_data;
  wire  ram_error__T_29_addr;
  wire  ram_error__T_29_mask;
  wire  ram_error__T_29_en;
  reg  value;
  reg [31:0] _RAND_5;
  reg  value_1;
  reg [31:0] _RAND_6;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_10;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_11;
  wire  _T_38;
  wire  _GEN_12;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_opcode = ram_opcode__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_source = ram_source__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign io_deq_bits_error = ram_error__T_43_data;
  assign ram_opcode__T_43_addr = value_1;
  assign ram_opcode__T_43_data = ram_opcode[ram_opcode__T_43_addr];
  assign ram_opcode__T_29_data = io_enq_bits_opcode;
  assign ram_opcode__T_29_addr = value;
  assign ram_opcode__T_29_mask = _T_25;
  assign ram_opcode__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_source__T_43_addr = value_1;
  assign ram_source__T_43_data = ram_source[ram_source__T_43_addr];
  assign ram_source__T_29_data = io_enq_bits_source;
  assign ram_source__T_29_addr = value;
  assign ram_source__T_29_mask = _T_25;
  assign ram_source__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign ram_error__T_43_addr = value_1;
  assign ram_error__T_43_data = ram_error[ram_error__T_43_addr];
  assign ram_error__T_29_data = io_enq_bits_error;
  assign ram_error__T_29_addr = value;
  assign ram_error__T_29_mask = _T_25;
  assign ram_error__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_10 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_11 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_12 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_3[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_error[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_29_en & ram_opcode__T_29_mask) begin
      ram_opcode[ram_opcode__T_29_addr] <= ram_opcode__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_source__T_29_en & ram_source__T_29_mask) begin
      ram_source[ram_source__T_29_addr] <= ram_source__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if(ram_error__T_29_en & ram_error__T_29_mask) begin
      ram_error[ram_error__T_29_addr] <= ram_error__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module TLBuffer_4(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input         io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output        io_in_0_d_bits_source,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output        io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input         io_out_0_d_bits_source,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [2:0] Queue_io_enq_bits_param;
  wire [3:0] Queue_io_enq_bits_size;
  wire  Queue_io_enq_bits_source;
  wire [31:0] Queue_io_enq_bits_address;
  wire [3:0] Queue_io_enq_bits_mask;
  wire [31:0] Queue_io_enq_bits_data;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [2:0] Queue_io_deq_bits_param;
  wire [3:0] Queue_io_deq_bits_size;
  wire  Queue_io_deq_bits_source;
  wire [31:0] Queue_io_deq_bits_address;
  wire [3:0] Queue_io_deq_bits_mask;
  wire [31:0] Queue_io_deq_bits_data;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [3:0] Queue_1_io_enq_bits_size;
  wire  Queue_1_io_enq_bits_source;
  wire [31:0] Queue_1_io_enq_bits_data;
  wire  Queue_1_io_enq_bits_error;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [3:0] Queue_1_io_deq_bits_size;
  wire  Queue_1_io_deq_bits_source;
  wire [31:0] Queue_1_io_deq_bits_data;
  wire  Queue_1_io_deq_bits_error;
  Queue_9 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_10 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_error(Queue_1_io_enq_bits_error),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_error(Queue_1_io_deq_bits_error)
  );
  assign io_in_0_a_ready = Queue_io_enq_ready;
  assign io_in_0_d_valid = Queue_1_io_deq_valid;
  assign io_in_0_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign io_in_0_d_bits_size = Queue_1_io_deq_bits_size;
  assign io_in_0_d_bits_source = Queue_1_io_deq_bits_source;
  assign io_in_0_d_bits_data = Queue_1_io_deq_bits_data;
  assign io_in_0_d_bits_error = Queue_1_io_deq_bits_error;
  assign io_out_0_a_valid = Queue_io_deq_valid;
  assign io_out_0_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign io_out_0_a_bits_param = Queue_io_deq_bits_param;
  assign io_out_0_a_bits_size = Queue_io_deq_bits_size;
  assign io_out_0_a_bits_source = Queue_io_deq_bits_source;
  assign io_out_0_a_bits_address = Queue_io_deq_bits_address;
  assign io_out_0_a_bits_mask = Queue_io_deq_bits_mask;
  assign io_out_0_a_bits_data = Queue_io_deq_bits_data;
  assign io_out_0_d_ready = Queue_1_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_a_valid;
  assign Queue_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Queue_io_enq_bits_param = io_in_0_a_bits_param;
  assign Queue_io_enq_bits_size = io_in_0_a_bits_size;
  assign Queue_io_enq_bits_source = io_in_0_a_bits_source;
  assign Queue_io_enq_bits_address = io_in_0_a_bits_address;
  assign Queue_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Queue_io_enq_bits_data = io_in_0_a_bits_data;
  assign Queue_io_deq_ready = io_out_0_a_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_out_0_d_valid;
  assign Queue_1_io_enq_bits_opcode = io_out_0_d_bits_opcode;
  assign Queue_1_io_enq_bits_size = io_out_0_d_bits_size;
  assign Queue_1_io_enq_bits_source = io_out_0_d_bits_source;
  assign Queue_1_io_enq_bits_data = io_out_0_d_bits_data;
  assign Queue_1_io_enq_bits_error = io_out_0_d_bits_error;
  assign Queue_1_io_deq_ready = io_in_0_d_ready;
endmodule
module IntXbar_1(
  input   io_in_0_0,
  output  io_out_0_0
);
  assign io_out_0_0 = io_in_0_0;
endmodule
module IntXbar_2(
  input   io_in_1_0,
  input   io_in_0_0,
  input   io_in_0_1,
  output  io_out_0_0,
  output  io_out_0_1,
  output  io_out_0_2
);
  assign io_out_0_0 = io_in_0_0;
  assign io_out_0_1 = io_in_0_1;
  assign io_out_0_2 = io_in_1_0;
endmodule
module IntXing(
  input   clock,
  input   io_in_0_0,
  input   io_in_0_1,
  output  io_out_0_0,
  output  io_out_0_1
);
  reg  _T_22_0;
  reg [31:0] _RAND_0;
  reg  _T_22_1;
  reg [31:0] _RAND_1;
  reg  _T_47_0;
  reg [31:0] _RAND_2;
  reg  _T_47_1;
  reg [31:0] _RAND_3;
  reg  _T_84_0;
  reg [31:0] _RAND_4;
  reg  _T_84_1;
  reg [31:0] _RAND_5;
  reg  _T_133_0;
  reg [31:0] _RAND_6;
  reg  _T_133_1;
  reg [31:0] _RAND_7;
  assign io_out_0_0 = _T_133_0;
  assign io_out_0_1 = _T_133_1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_22_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_22_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_47_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_47_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_84_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_84_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_133_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_133_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_22_0 <= io_in_0_0;
    _T_22_1 <= io_in_0_1;
    _T_47_0 <= _T_22_0;
    _T_47_1 <= _T_22_1;
    _T_84_0 <= _T_47_0;
    _T_84_1 <= _T_47_1;
    _T_133_0 <= _T_84_0;
    _T_133_1 <= _T_84_1;
  end
endmodule
module Queue_11(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
  reg [63:0] ram_data [0:0];
  reg [63:0] _RAND_0;
  wire [63:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [63:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg [7:0] ram_strb [0:0];
  reg [31:0] _RAND_1;
  wire [7:0] ram_strb__T_35_data;
  wire  ram_strb__T_35_addr;
  wire [7:0] ram_strb__T_26_data;
  wire  ram_strb__T_26_addr;
  wire  ram_strb__T_26_mask;
  wire  ram_strb__T_26_en;
  reg  ram_last [0:0];
  reg [31:0] _RAND_2;
  wire  ram_last__T_35_data;
  wire  ram_last__T_35_addr;
  wire  ram_last__T_26_data;
  wire  ram_last__T_26_addr;
  wire  ram_last__T_26_mask;
  wire  ram_last__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_6;
  wire  _T_31;
  wire  _GEN_7;
  wire  _GEN_8;
  wire [63:0] _GEN_9;
  wire [7:0] _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_7;
  assign io_deq_bits_data = _GEN_9;
  assign io_deq_bits_strb = _GEN_10;
  assign io_deq_bits_last = _GEN_11;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _GEN_13;
  assign ram_data__T_26_en = _GEN_13;
  assign ram_strb__T_35_addr = 1'h0;
  assign ram_strb__T_35_data = ram_strb[ram_strb__T_35_addr];
  assign ram_strb__T_26_data = io_enq_bits_strb;
  assign ram_strb__T_26_addr = 1'h0;
  assign ram_strb__T_26_mask = _GEN_13;
  assign ram_strb__T_26_en = _GEN_13;
  assign ram_last__T_35_addr = 1'h0;
  assign ram_last__T_35_data = ram_last[ram_last__T_35_addr];
  assign ram_last__T_26_data = io_enq_bits_last;
  assign ram_last__T_26_addr = 1'h0;
  assign ram_last__T_26_mask = _GEN_13;
  assign ram_last__T_26_en = _GEN_13;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_13 != _GEN_12;
  assign _GEN_6 = _T_29 ? _GEN_13 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_7 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_8 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_9 = _T_18 ? io_enq_bits_data : ram_data__T_35_data;
  assign _GEN_10 = _T_18 ? io_enq_bits_strb : ram_strb__T_35_data;
  assign _GEN_11 = _T_18 ? io_enq_bits_last : ram_last__T_35_data;
  assign _GEN_12 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_13 = _T_18 ? _GEN_8 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if(ram_strb__T_26_en & ram_strb__T_26_mask) begin
      ram_strb[ram_strb__T_26_addr] <= ram_strb__T_26_data;
    end
    if(ram_last__T_26_en & ram_last__T_26_mask) begin
      ram_last[ram_last__T_26_addr] <= ram_last__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_12(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [1:0]  io_enq_bits_id,
  input  [30:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [11:0] io_enq_bits_user,
  input         io_enq_bits_wen,
  input         io_deq_ready,
  output        io_deq_valid,
  output [1:0]  io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [11:0] io_deq_bits_user,
  output        io_deq_bits_wen
);
  reg [1:0] ram_id [0:0];
  reg [31:0] _RAND_0;
  wire [1:0] ram_id__T_35_data;
  wire  ram_id__T_35_addr;
  wire [1:0] ram_id__T_26_data;
  wire  ram_id__T_26_addr;
  wire  ram_id__T_26_mask;
  wire  ram_id__T_26_en;
  reg [30:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [30:0] ram_addr__T_35_data;
  wire  ram_addr__T_35_addr;
  wire [30:0] ram_addr__T_26_data;
  wire  ram_addr__T_26_addr;
  wire  ram_addr__T_26_mask;
  wire  ram_addr__T_26_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_35_data;
  wire  ram_len__T_35_addr;
  wire [7:0] ram_len__T_26_data;
  wire  ram_len__T_26_addr;
  wire  ram_len__T_26_mask;
  wire  ram_len__T_26_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [2:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_35_data;
  wire  ram_burst__T_35_addr;
  wire [1:0] ram_burst__T_26_data;
  wire  ram_burst__T_26_addr;
  wire  ram_burst__T_26_mask;
  wire  ram_burst__T_26_en;
  reg [11:0] ram_user [0:0];
  reg [31:0] _RAND_5;
  wire [11:0] ram_user__T_35_data;
  wire  ram_user__T_35_addr;
  wire [11:0] ram_user__T_26_data;
  wire  ram_user__T_26_addr;
  wire  ram_user__T_26_mask;
  wire  ram_user__T_26_en;
  reg  ram_wen [0:0];
  reg [31:0] _RAND_6;
  wire  ram_wen__T_35_data;
  wire  ram_wen__T_35_addr;
  wire  ram_wen__T_26_data;
  wire  ram_wen__T_26_addr;
  wire  ram_wen__T_26_mask;
  wire  ram_wen__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_14;
  wire  _T_31;
  wire  _GEN_15;
  wire  _GEN_16;
  wire [1:0] _GEN_17;
  wire [30:0] _GEN_18;
  wire [7:0] _GEN_19;
  wire [2:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [11:0] _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_15;
  assign io_deq_bits_id = _GEN_17;
  assign io_deq_bits_addr = _GEN_18;
  assign io_deq_bits_len = _GEN_19;
  assign io_deq_bits_size = _GEN_20;
  assign io_deq_bits_burst = _GEN_21;
  assign io_deq_bits_user = _GEN_26;
  assign io_deq_bits_wen = _GEN_27;
  assign ram_id__T_35_addr = 1'h0;
  assign ram_id__T_35_data = ram_id[ram_id__T_35_addr];
  assign ram_id__T_26_data = io_enq_bits_id;
  assign ram_id__T_26_addr = 1'h0;
  assign ram_id__T_26_mask = _GEN_29;
  assign ram_id__T_26_en = _GEN_29;
  assign ram_addr__T_35_addr = 1'h0;
  assign ram_addr__T_35_data = ram_addr[ram_addr__T_35_addr];
  assign ram_addr__T_26_data = io_enq_bits_addr;
  assign ram_addr__T_26_addr = 1'h0;
  assign ram_addr__T_26_mask = _GEN_29;
  assign ram_addr__T_26_en = _GEN_29;
  assign ram_len__T_35_addr = 1'h0;
  assign ram_len__T_35_data = ram_len[ram_len__T_35_addr];
  assign ram_len__T_26_data = io_enq_bits_len;
  assign ram_len__T_26_addr = 1'h0;
  assign ram_len__T_26_mask = _GEN_29;
  assign ram_len__T_26_en = _GEN_29;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_29;
  assign ram_size__T_26_en = _GEN_29;
  assign ram_burst__T_35_addr = 1'h0;
  assign ram_burst__T_35_data = ram_burst[ram_burst__T_35_addr];
  assign ram_burst__T_26_data = io_enq_bits_burst;
  assign ram_burst__T_26_addr = 1'h0;
  assign ram_burst__T_26_mask = _GEN_29;
  assign ram_burst__T_26_en = _GEN_29;
  assign ram_user__T_35_addr = 1'h0;
  assign ram_user__T_35_data = ram_user[ram_user__T_35_addr];
  assign ram_user__T_26_data = io_enq_bits_user;
  assign ram_user__T_26_addr = 1'h0;
  assign ram_user__T_26_mask = _GEN_29;
  assign ram_user__T_26_en = _GEN_29;
  assign ram_wen__T_35_addr = 1'h0;
  assign ram_wen__T_35_data = ram_wen[ram_wen__T_35_addr];
  assign ram_wen__T_26_data = io_enq_bits_wen;
  assign ram_wen__T_26_addr = 1'h0;
  assign ram_wen__T_26_mask = _GEN_29;
  assign ram_wen__T_26_en = _GEN_29;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_29 != _GEN_28;
  assign _GEN_14 = _T_29 ? _GEN_29 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_15 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_16 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_17 = _T_18 ? io_enq_bits_id : ram_id__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_addr : ram_addr__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_len : ram_len__T_35_data;
  assign _GEN_20 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_21 = _T_18 ? io_enq_bits_burst : ram_burst__T_35_data;
  assign _GEN_26 = _T_18 ? io_enq_bits_user : ram_user__T_35_data;
  assign _GEN_27 = _T_18 ? io_enq_bits_wen : ram_wen__T_35_data;
  assign _GEN_28 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_29 = _T_18 ? _GEN_16 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = _RAND_5[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_wen[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_26_en & ram_id__T_26_mask) begin
      ram_id[ram_id__T_26_addr] <= ram_id__T_26_data;
    end
    if(ram_addr__T_26_en & ram_addr__T_26_mask) begin
      ram_addr[ram_addr__T_26_addr] <= ram_addr__T_26_data;
    end
    if(ram_len__T_26_en & ram_len__T_26_mask) begin
      ram_len[ram_len__T_26_addr] <= ram_len__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_burst__T_26_en & ram_burst__T_26_mask) begin
      ram_burst[ram_burst__T_26_addr] <= ram_burst__T_26_data;
    end
    if(ram_user__T_26_en & ram_user__T_26_mask) begin
      ram_user[ram_user__T_26_addr] <= ram_user__T_26_data;
    end
    if(ram_wen__T_26_en & ram_wen__T_26_mask) begin
      ram_wen[ram_wen__T_26_addr] <= ram_wen__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module TLToAXI4(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [3:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input  [30:0] io_in_0_a_bits_address,
  input  [7:0]  io_in_0_a_bits_mask,
  input  [63:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [3:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [63:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [1:0]  io_out_0_aw_bits_id,
  output [30:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [1:0]  io_out_0_aw_bits_burst,
  output [11:0] io_out_0_aw_bits_user,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [1:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input  [11:0] io_out_0_b_bits_user,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [1:0]  io_out_0_ar_bits_id,
  output [30:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [1:0]  io_out_0_ar_bits_burst,
  output [11:0] io_out_0_ar_bits_user,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [1:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input  [11:0] io_out_0_r_bits_user,
  input         io_out_0_r_bits_last
);
  wire  _T_197;
  wire  _T_199;
  wire  _T_200;
  wire [22:0] _T_203;
  wire [7:0] _T_204;
  wire [7:0] _T_205;
  wire [4:0] _T_206;
  wire [4:0] _T_211;
  reg [4:0] _T_214;
  reg [31:0] _RAND_0;
  wire [5:0] _T_216;
  wire [5:0] _T_217;
  wire [4:0] _T_218;
  wire  _T_220;
  wire  _T_222;
  wire  _T_224;
  wire  _T_225;
  wire [4:0] _T_229;
  wire [4:0] _GEN_4;
  wire [8:0] _GEN_43;
  wire [8:0] _T_241;
  wire [8:0] _GEN_44;
  wire [8:0] _T_242;
  wire [4:0] _T_243;
  wire [3:0] _T_244;
  wire [4:0] _T_245;
  wire [3:0] _T_246;
  wire  _T_252_ready;
  wire [2:0] _T_252_bits_size;
  wire [11:0] _T_252_bits_user;
  wire  _T_256_ready;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [63:0] Queue_io_enq_bits_data;
  wire [7:0] Queue_io_enq_bits_strb;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [63:0] Queue_io_deq_bits_data;
  wire [7:0] Queue_io_deq_bits_strb;
  wire  Queue_io_deq_bits_last;
  wire  _T_265_valid;
  wire [63:0] _T_265_bits_data;
  wire [7:0] _T_265_bits_strb;
  wire  _T_265_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [1:0] Queue_1_io_enq_bits_id;
  wire [30:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [1:0] Queue_1_io_enq_bits_burst;
  wire [11:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_enq_bits_wen;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [1:0] Queue_1_io_deq_bits_id;
  wire [30:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire [11:0] Queue_1_io_deq_bits_user;
  wire  Queue_1_io_deq_bits_wen;
  wire  _T_274_valid;
  wire [1:0] _T_274_bits_id;
  wire [30:0] _T_274_bits_addr;
  wire [7:0] _T_274_bits_len;
  wire [2:0] _T_274_bits_size;
  wire [1:0] _T_274_bits_burst;
  wire [11:0] _T_274_bits_user;
  wire  _T_274_bits_wen;
  wire  _T_279;
  wire  _T_280;
  wire  _T_281;
  wire  _T_282;
  reg  _T_286;
  reg [31:0] _RAND_1;
  wire  _T_289;
  wire  _GEN_5;
  wire [1:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [1:0] _GEN_16;
  wire [1:0] _GEN_17;
  wire [1:0] _GEN_18;
  wire [1:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [1:0] _GEN_22;
  wire [25:0] _T_293;
  wire [10:0] _T_294;
  wire [10:0] _T_295;
  wire [7:0] _T_296;
  wire  _T_297;
  wire [3:0] _T_298;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire  _T_306;
  wire  _T_307;
  wire  _T_308;
  wire  _T_309;
  wire  _T_310;
  wire  _T_313;
  wire  _T_315;
  wire  _T_316;
  wire  _T_318;
  wire  _T_319;
  wire  _T_323;
  wire  _T_325;
  reg  _T_328;
  reg [31:0] _RAND_2;
  wire  _T_329;
  wire  _T_331;
  wire  _GEN_40;
  wire  _T_332;
  wire  _T_334;
  wire  _T_335;
  wire  _T_336;
  wire  _T_338;
  wire  _T_340;
  wire [2:0] _T_353_opcode;
  wire [3:0] _T_353_size;
  wire [4:0] _T_353_source;
  wire  _T_353_error;
  wire [3:0] _T_356;
  wire  _T_360;
  wire  _T_361;
  wire [1:0] _T_362;
  wire [3:0] _T_365;
  wire  _T_369;
  wire  _T_370;
  wire  _T_372;
  reg [3:0] _T_375;
  reg [31:0] _RAND_3;
  reg  _T_377;
  reg [31:0] _RAND_4;
  wire  _T_379;
  wire  _T_380;
  wire  _T_381;
  wire  _T_382;
  wire  _T_383;
  wire  _T_384;
  wire [3:0] _GEN_45;
  wire [4:0] _T_385;
  wire [3:0] _T_386;
  wire [3:0] _GEN_46;
  wire [4:0] _T_387;
  wire [4:0] _T_388;
  wire [3:0] _T_389;
  wire  _T_391;
  wire  _T_393;
  wire  _T_394;
  wire  _T_395;
  wire  _T_397;
  wire  _T_399;
  wire  _T_401;
  wire  _T_402;
  wire  _T_403;
  wire  _T_405;
  wire  _GEN_41;
  wire  _T_407;
  wire  _T_408;
  wire  _T_409;
  reg [3:0] _T_412;
  reg [31:0] _RAND_5;
  reg  _T_414;
  reg [31:0] _RAND_6;
  wire  _T_416;
  wire  _T_418;
  wire  _T_419;
  wire  _T_421;
  wire [3:0] _GEN_47;
  wire [4:0] _T_422;
  wire [3:0] _T_423;
  wire [3:0] _GEN_48;
  wire [4:0] _T_424;
  wire [4:0] _T_425;
  wire [3:0] _T_426;
  wire  _T_428;
  wire  _T_430;
  wire  _T_431;
  wire  _T_432;
  wire  _T_434;
  wire  _T_436;
  wire  _T_438;
  wire  _T_439;
  wire  _T_440;
  wire  _T_442;
  wire  _GEN_42;
  wire  _T_444;
  wire  _T_445;
  wire  _T_446;
  Queue_11 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_strb(Queue_io_enq_bits_strb),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_strb(Queue_io_deq_bits_strb),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_12 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_wen(Queue_1_io_enq_bits_wen),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_wen(Queue_1_io_deq_bits_wen)
  );
  assign io_in_0_a_ready = _T_310;
  assign io_in_0_d_valid = _T_336;
  assign io_in_0_d_bits_opcode = _T_353_opcode;
  assign io_in_0_d_bits_param = 2'h0;
  assign io_in_0_d_bits_size = _T_353_size;
  assign io_in_0_d_bits_source = _T_353_source;
  assign io_in_0_d_bits_sink = 1'h0;
  assign io_in_0_d_bits_data = io_out_0_r_bits_data;
  assign io_in_0_d_bits_error = _T_353_error;
  assign io_out_0_aw_valid = _T_281;
  assign io_out_0_aw_bits_id = _T_274_bits_id;
  assign io_out_0_aw_bits_addr = _T_274_bits_addr;
  assign io_out_0_aw_bits_len = _T_274_bits_len;
  assign io_out_0_aw_bits_size = _T_274_bits_size;
  assign io_out_0_aw_bits_burst = _T_274_bits_burst;
  assign io_out_0_aw_bits_user = _T_274_bits_user;
  assign io_out_0_w_valid = _T_265_valid;
  assign io_out_0_w_bits_data = _T_265_bits_data;
  assign io_out_0_w_bits_strb = _T_265_bits_strb;
  assign io_out_0_w_bits_last = _T_265_bits_last;
  assign io_out_0_b_ready = _T_335;
  assign io_out_0_ar_valid = _T_280;
  assign io_out_0_ar_bits_id = _T_274_bits_id;
  assign io_out_0_ar_bits_addr = _T_274_bits_addr;
  assign io_out_0_ar_bits_len = _T_274_bits_len;
  assign io_out_0_ar_bits_size = _T_274_bits_size;
  assign io_out_0_ar_bits_burst = _T_274_bits_burst;
  assign io_out_0_ar_bits_user = _T_274_bits_user;
  assign io_out_0_r_ready = io_in_0_d_ready;
  assign _T_197 = io_in_0_a_bits_opcode[2];
  assign _T_199 = _T_197 == 1'h0;
  assign _T_200 = io_in_0_a_ready & io_in_0_a_valid;
  assign _T_203 = 23'hff << io_in_0_a_bits_size;
  assign _T_204 = _T_203[7:0];
  assign _T_205 = ~ _T_204;
  assign _T_206 = _T_205[7:3];
  assign _T_211 = _T_199 ? _T_206 : 5'h0;
  assign _T_216 = _T_214 - 5'h1;
  assign _T_217 = $unsigned(_T_216);
  assign _T_218 = _T_217[4:0];
  assign _T_220 = _T_214 == 5'h0;
  assign _T_222 = _T_214 == 5'h1;
  assign _T_224 = _T_211 == 5'h0;
  assign _T_225 = _T_222 | _T_224;
  assign _T_229 = _T_220 ? _T_211 : _T_218;
  assign _GEN_4 = _T_200 ? _T_229 : _T_214;
  assign _GEN_43 = {{5'd0}, io_in_0_a_bits_size};
  assign _T_241 = _GEN_43 << 5;
  assign _GEN_44 = {{4'd0}, io_in_0_a_bits_source};
  assign _T_242 = _GEN_44 | _T_241;
  assign _T_243 = io_out_0_r_bits_user[4:0];
  assign _T_244 = io_out_0_r_bits_user[8:5];
  assign _T_245 = io_out_0_b_bits_user[4:0];
  assign _T_246 = io_out_0_b_bits_user[8:5];
  assign _T_252_ready = Queue_1_io_enq_ready;
  assign _T_252_bits_size = _T_298[2:0];
  assign _T_252_bits_user = {{3'd0}, _T_242};
  assign _T_256_ready = Queue_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_325;
  assign Queue_io_enq_bits_data = io_in_0_a_bits_data;
  assign Queue_io_enq_bits_strb = io_in_0_a_bits_mask;
  assign Queue_io_enq_bits_last = _T_225;
  assign Queue_io_deq_ready = io_out_0_w_ready;
  assign _T_265_valid = Queue_io_deq_valid;
  assign _T_265_bits_data = Queue_io_deq_bits_data;
  assign _T_265_bits_strb = Queue_io_deq_bits_strb;
  assign _T_265_bits_last = Queue_io_deq_bits_last;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_319;
  assign Queue_1_io_enq_bits_id = _GEN_22;
  assign Queue_1_io_enq_bits_addr = io_in_0_a_bits_address;
  assign Queue_1_io_enq_bits_len = _T_296;
  assign Queue_1_io_enq_bits_size = _T_252_bits_size;
  assign Queue_1_io_enq_bits_burst = 2'h1;
  assign Queue_1_io_enq_bits_user = _T_252_bits_user;
  assign Queue_1_io_enq_bits_wen = _T_199;
  assign Queue_1_io_deq_ready = _T_282;
  assign _T_274_valid = Queue_1_io_deq_valid;
  assign _T_274_bits_id = Queue_1_io_deq_bits_id;
  assign _T_274_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_274_bits_len = Queue_1_io_deq_bits_len;
  assign _T_274_bits_size = Queue_1_io_deq_bits_size;
  assign _T_274_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_274_bits_user = Queue_1_io_deq_bits_user;
  assign _T_274_bits_wen = Queue_1_io_deq_bits_wen;
  assign _T_279 = _T_274_bits_wen == 1'h0;
  assign _T_280 = _T_274_valid & _T_279;
  assign _T_281 = _T_274_valid & _T_274_bits_wen;
  assign _T_282 = _T_274_bits_wen ? io_out_0_aw_ready : io_out_0_ar_ready;
  assign _T_289 = _T_225 == 1'h0;
  assign _GEN_5 = _T_200 ? _T_289 : _T_286;
  assign _GEN_13 = 5'h8 == io_in_0_a_bits_source ? 2'h3 : 2'h2;
  assign _GEN_14 = 5'h9 == io_in_0_a_bits_source ? 2'h3 : _GEN_13;
  assign _GEN_15 = 5'ha == io_in_0_a_bits_source ? 2'h3 : _GEN_14;
  assign _GEN_16 = 5'hb == io_in_0_a_bits_source ? 2'h3 : _GEN_15;
  assign _GEN_17 = 5'hc == io_in_0_a_bits_source ? 2'h3 : _GEN_16;
  assign _GEN_18 = 5'hd == io_in_0_a_bits_source ? 2'h3 : _GEN_17;
  assign _GEN_19 = 5'he == io_in_0_a_bits_source ? 2'h3 : _GEN_18;
  assign _GEN_20 = 5'hf == io_in_0_a_bits_source ? 2'h3 : _GEN_19;
  assign _GEN_21 = 5'h10 == io_in_0_a_bits_source ? 2'h0 : _GEN_20;
  assign _GEN_22 = 5'h11 == io_in_0_a_bits_source ? 2'h1 : _GEN_21;
  assign _T_293 = 26'h7ff << io_in_0_a_bits_size;
  assign _T_294 = _T_293[10:0];
  assign _T_295 = ~ _T_294;
  assign _T_296 = _T_295[10:3];
  assign _T_297 = io_in_0_a_bits_size >= 4'h3;
  assign _T_298 = _T_297 ? 4'h3 : io_in_0_a_bits_size;
  assign _GEN_30 = 5'h8 == io_in_0_a_bits_source ? _T_446 : _T_409;
  assign _GEN_31 = 5'h9 == io_in_0_a_bits_source ? _T_446 : _GEN_30;
  assign _GEN_32 = 5'ha == io_in_0_a_bits_source ? _T_446 : _GEN_31;
  assign _GEN_33 = 5'hb == io_in_0_a_bits_source ? _T_446 : _GEN_32;
  assign _GEN_34 = 5'hc == io_in_0_a_bits_source ? _T_446 : _GEN_33;
  assign _GEN_35 = 5'hd == io_in_0_a_bits_source ? _T_446 : _GEN_34;
  assign _GEN_36 = 5'he == io_in_0_a_bits_source ? _T_446 : _GEN_35;
  assign _GEN_37 = 5'hf == io_in_0_a_bits_source ? _T_446 : _GEN_36;
  assign _GEN_38 = 5'h10 == io_in_0_a_bits_source ? 1'h0 : _GEN_37;
  assign _GEN_39 = 5'h11 == io_in_0_a_bits_source ? 1'h0 : _GEN_38;
  assign _T_306 = _GEN_39 == 1'h0;
  assign _T_307 = _T_286 | _T_252_ready;
  assign _T_308 = _T_307 & _T_256_ready;
  assign _T_309 = _T_199 ? _T_308 : _T_252_ready;
  assign _T_310 = _T_306 & _T_309;
  assign _T_313 = _T_306 & io_in_0_a_valid;
  assign _T_315 = _T_286 == 1'h0;
  assign _T_316 = _T_315 & _T_256_ready;
  assign _T_318 = _T_199 ? _T_316 : 1'h1;
  assign _T_319 = _T_313 & _T_318;
  assign _T_323 = _T_313 & _T_199;
  assign _T_325 = _T_323 & _T_307;
  assign _T_329 = io_out_0_r_ready & io_out_0_r_valid;
  assign _T_331 = io_out_0_r_bits_last == 1'h0;
  assign _GEN_40 = _T_329 ? _T_331 : _T_328;
  assign _T_332 = io_out_0_r_valid | _T_328;
  assign _T_334 = _T_332 == 1'h0;
  assign _T_335 = io_in_0_d_ready & _T_334;
  assign _T_336 = _T_332 ? io_out_0_r_valid : io_out_0_b_valid;
  assign _T_338 = io_out_0_r_bits_resp != 2'h0;
  assign _T_340 = io_out_0_b_bits_resp != 2'h0;
  assign _T_353_opcode = _T_332 ? 3'h1 : 3'h0;
  assign _T_353_size = _T_332 ? _T_244 : _T_246;
  assign _T_353_source = _T_332 ? _T_243 : _T_245;
  assign _T_353_error = _T_332 ? _T_338 : _T_340;
  assign _T_356 = 4'h1 << _GEN_22;
  assign _T_360 = _T_356[2];
  assign _T_361 = _T_356[3];
  assign _T_362 = _T_332 ? io_out_0_r_bits_id : io_out_0_b_bits_id;
  assign _T_365 = 4'h1 << _T_362;
  assign _T_369 = _T_365[2];
  assign _T_370 = _T_365[3];
  assign _T_372 = _T_332 ? io_out_0_r_bits_last : 1'h1;
  assign _T_379 = _T_375 == 4'h0;
  assign _T_380 = _T_252_ready & _T_319;
  assign _T_381 = _T_360 & _T_380;
  assign _T_382 = _T_369 & _T_372;
  assign _T_383 = io_in_0_d_ready & io_in_0_d_valid;
  assign _T_384 = _T_382 & _T_383;
  assign _GEN_45 = {{3'd0}, _T_381};
  assign _T_385 = _T_375 + _GEN_45;
  assign _T_386 = _T_385[3:0];
  assign _GEN_46 = {{3'd0}, _T_384};
  assign _T_387 = _T_386 - _GEN_46;
  assign _T_388 = $unsigned(_T_387);
  assign _T_389 = _T_388[3:0];
  assign _T_391 = _T_384 == 1'h0;
  assign _T_393 = _T_375 != 4'h0;
  assign _T_394 = _T_391 | _T_393;
  assign _T_395 = _T_394 | reset;
  assign _T_397 = _T_395 == 1'h0;
  assign _T_399 = _T_381 == 1'h0;
  assign _T_401 = _T_375 != 4'h8;
  assign _T_402 = _T_399 | _T_401;
  assign _T_403 = _T_402 | reset;
  assign _T_405 = _T_403 == 1'h0;
  assign _GEN_41 = _T_381 ? _T_199 : _T_377;
  assign _T_407 = _T_379 == 1'h0;
  assign _T_408 = _T_377 != _T_199;
  assign _T_409 = _T_407 & _T_408;
  assign _T_416 = _T_412 == 4'h0;
  assign _T_418 = _T_361 & _T_380;
  assign _T_419 = _T_370 & _T_372;
  assign _T_421 = _T_419 & _T_383;
  assign _GEN_47 = {{3'd0}, _T_418};
  assign _T_422 = _T_412 + _GEN_47;
  assign _T_423 = _T_422[3:0];
  assign _GEN_48 = {{3'd0}, _T_421};
  assign _T_424 = _T_423 - _GEN_48;
  assign _T_425 = $unsigned(_T_424);
  assign _T_426 = _T_425[3:0];
  assign _T_428 = _T_421 == 1'h0;
  assign _T_430 = _T_412 != 4'h0;
  assign _T_431 = _T_428 | _T_430;
  assign _T_432 = _T_431 | reset;
  assign _T_434 = _T_432 == 1'h0;
  assign _T_436 = _T_418 == 1'h0;
  assign _T_438 = _T_412 != 4'h8;
  assign _T_439 = _T_436 | _T_438;
  assign _T_440 = _T_439 | reset;
  assign _T_442 = _T_440 == 1'h0;
  assign _GEN_42 = _T_418 ? _T_199 : _T_414;
  assign _T_444 = _T_416 == 1'h0;
  assign _T_445 = _T_414 != _T_199;
  assign _T_446 = _T_444 & _T_445;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_214 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_286 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_328 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_375 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_377 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_412 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_414 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_214 <= 5'h0;
    end else begin
      if (_T_200) begin
        if (_T_220) begin
          if (_T_199) begin
            _T_214 <= _T_206;
          end else begin
            _T_214 <= 5'h0;
          end
        end else begin
          _T_214 <= _T_218;
        end
      end
    end
    if (reset) begin
      _T_286 <= 1'h0;
    end else begin
      if (_T_200) begin
        _T_286 <= _T_289;
      end
    end
    if (reset) begin
      _T_328 <= 1'h0;
    end else begin
      if (_T_329) begin
        _T_328 <= _T_331;
      end
    end
    if (reset) begin
      _T_375 <= 4'h0;
    end else begin
      _T_375 <= _T_389;
    end
    if (_T_381) begin
      _T_377 <= _T_199;
    end
    if (reset) begin
      _T_412 <= 4'h0;
    end else begin
      _T_412 <= _T_426;
    end
    if (_T_418) begin
      _T_414 <= _T_199;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:112 assert (a_source  < UInt(BigInt(1) << sourceBits))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:113 assert (a_size    < UInt(BigInt(1) << sizeBits))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_397) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:206 assert (!dec || count =/= UInt(0))     // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_397) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_405) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:207 assert (!inc || count =/= UInt(n.get)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_405) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_434) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:206 assert (!dec || count =/= UInt(0))     // underflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_434) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_442) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:207 assert (!inc || count =/= UInt(n.get)) // overflow\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_442) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4IdIndexer(
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [1:0]  io_in_0_aw_bits_id,
  input  [30:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  input  [11:0] io_in_0_aw_bits_user,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [1:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output [11:0] io_in_0_b_bits_user,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [1:0]  io_in_0_ar_bits_id,
  input  [30:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input  [11:0] io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [1:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output [11:0] io_in_0_r_bits_user,
  output        io_in_0_r_bits_last,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [3:0]  io_out_0_aw_bits_id,
  output [30:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [1:0]  io_out_0_aw_bits_burst,
  output [11:0] io_out_0_aw_bits_user,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [3:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input  [11:0] io_out_0_b_bits_user,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [3:0]  io_out_0_ar_bits_id,
  output [30:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [1:0]  io_out_0_ar_bits_burst,
  output [11:0] io_out_0_ar_bits_user,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [3:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input  [11:0] io_out_0_r_bits_user,
  input         io_out_0_r_bits_last
);
  assign io_in_0_aw_ready = io_out_0_aw_ready;
  assign io_in_0_w_ready = io_out_0_w_ready;
  assign io_in_0_b_valid = io_out_0_b_valid;
  assign io_in_0_b_bits_id = io_out_0_b_bits_id[1:0];
  assign io_in_0_b_bits_resp = io_out_0_b_bits_resp;
  assign io_in_0_b_bits_user = io_out_0_b_bits_user;
  assign io_in_0_ar_ready = io_out_0_ar_ready;
  assign io_in_0_r_valid = io_out_0_r_valid;
  assign io_in_0_r_bits_id = io_out_0_r_bits_id[1:0];
  assign io_in_0_r_bits_data = io_out_0_r_bits_data;
  assign io_in_0_r_bits_resp = io_out_0_r_bits_resp;
  assign io_in_0_r_bits_user = io_out_0_r_bits_user;
  assign io_in_0_r_bits_last = io_out_0_r_bits_last;
  assign io_out_0_aw_valid = io_in_0_aw_valid;
  assign io_out_0_aw_bits_id = {{2'd0}, io_in_0_aw_bits_id};
  assign io_out_0_aw_bits_addr = io_in_0_aw_bits_addr;
  assign io_out_0_aw_bits_len = io_in_0_aw_bits_len;
  assign io_out_0_aw_bits_size = io_in_0_aw_bits_size;
  assign io_out_0_aw_bits_burst = io_in_0_aw_bits_burst;
  assign io_out_0_aw_bits_user = io_in_0_aw_bits_user;
  assign io_out_0_w_valid = io_in_0_w_valid;
  assign io_out_0_w_bits_data = io_in_0_w_bits_data;
  assign io_out_0_w_bits_strb = io_in_0_w_bits_strb;
  assign io_out_0_w_bits_last = io_in_0_w_bits_last;
  assign io_out_0_b_ready = io_in_0_b_ready;
  assign io_out_0_ar_valid = io_in_0_ar_valid;
  assign io_out_0_ar_bits_id = {{2'd0}, io_in_0_ar_bits_id};
  assign io_out_0_ar_bits_addr = io_in_0_ar_bits_addr;
  assign io_out_0_ar_bits_len = io_in_0_ar_bits_len;
  assign io_out_0_ar_bits_size = io_in_0_ar_bits_size;
  assign io_out_0_ar_bits_burst = io_in_0_ar_bits_burst;
  assign io_out_0_ar_bits_user = io_in_0_ar_bits_user;
  assign io_out_0_r_ready = io_in_0_r_ready;
endmodule
module Queue_13(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input  [11:0] io_enq_bits_user,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output [11:0] io_deq_bits_user,
  output        io_deq_bits_last
);
  reg [3:0] ram_id [0:7];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire [2:0] ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire [2:0] ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [63:0] ram_data [0:7];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_43_data;
  wire [2:0] ram_data__T_43_addr;
  wire [63:0] ram_data__T_29_data;
  wire [2:0] ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg [1:0] ram_resp [0:7];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_43_data;
  wire [2:0] ram_resp__T_43_addr;
  wire [1:0] ram_resp__T_29_data;
  wire [2:0] ram_resp__T_29_addr;
  wire  ram_resp__T_29_mask;
  wire  ram_resp__T_29_en;
  reg [11:0] ram_user [0:7];
  reg [31:0] _RAND_3;
  wire [11:0] ram_user__T_43_data;
  wire [2:0] ram_user__T_43_addr;
  wire [11:0] ram_user__T_29_data;
  wire [2:0] ram_user__T_29_addr;
  wire  ram_user__T_29_mask;
  wire  ram_user__T_29_en;
  reg  ram_last [0:7];
  reg [31:0] _RAND_4;
  wire  ram_last__T_43_data;
  wire [2:0] ram_last__T_43_addr;
  wire  ram_last__T_29_data;
  wire [2:0] ram_last__T_29_addr;
  wire  ram_last__T_29_mask;
  wire  ram_last__T_29_en;
  reg [2:0] value;
  reg [31:0] _RAND_5;
  reg [2:0] value_1;
  reg [31:0] _RAND_6;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [3:0] _T_32;
  wire [2:0] _T_33;
  wire [2:0] _GEN_8;
  wire [3:0] _T_36;
  wire [2:0] _T_37;
  wire [2:0] _GEN_9;
  wire  _T_38;
  wire  _GEN_10;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign io_deq_bits_resp = ram_resp__T_43_data;
  assign io_deq_bits_user = ram_user__T_43_data;
  assign io_deq_bits_last = ram_last__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign ram_resp__T_43_addr = value_1;
  assign ram_resp__T_43_data = ram_resp[ram_resp__T_43_addr];
  assign ram_resp__T_29_data = io_enq_bits_resp;
  assign ram_resp__T_29_addr = value;
  assign ram_resp__T_29_mask = _T_25;
  assign ram_resp__T_29_en = _T_25;
  assign ram_user__T_43_addr = value_1;
  assign ram_user__T_43_data = ram_user[ram_user__T_43_addr];
  assign ram_user__T_29_data = io_enq_bits_user;
  assign ram_user__T_29_addr = value;
  assign ram_user__T_29_mask = _T_25;
  assign ram_user__T_29_en = _T_25;
  assign ram_last__T_43_addr = value_1;
  assign ram_last__T_43_data = ram_last[ram_last__T_43_addr];
  assign ram_last__T_29_data = io_enq_bits_last;
  assign ram_last__T_29_addr = value;
  assign ram_last__T_29_mask = _T_25;
  assign ram_last__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 3'h1;
  assign _T_33 = _T_32[2:0];
  assign _GEN_8 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 3'h1;
  assign _T_37 = _T_36[2:0];
  assign _GEN_9 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_10 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_user[initvar] = _RAND_3[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram_last[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value_1 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if(ram_resp__T_29_en & ram_resp__T_29_mask) begin
      ram_resp[ram_resp__T_29_addr] <= ram_resp__T_29_data;
    end
    if(ram_user__T_29_en & ram_user__T_29_mask) begin
      ram_user[ram_user__T_29_addr] <= ram_user__T_29_data;
    end
    if(ram_last__T_29_en & ram_last__T_29_mask) begin
      ram_last[ram_last__T_29_addr] <= ram_last__T_29_data;
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module AXI4Deinterleaver(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [3:0]  io_in_0_aw_bits_id,
  input  [30:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  input  [11:0] io_in_0_aw_bits_user,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [3:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output [11:0] io_in_0_b_bits_user,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [3:0]  io_in_0_ar_bits_id,
  input  [30:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input  [11:0] io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [3:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output [11:0] io_in_0_r_bits_user,
  output        io_in_0_r_bits_last,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [3:0]  io_out_0_aw_bits_id,
  output [30:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [1:0]  io_out_0_aw_bits_burst,
  output [11:0] io_out_0_aw_bits_user,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [3:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input  [11:0] io_out_0_b_bits_user,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [3:0]  io_out_0_ar_bits_id,
  output [30:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [1:0]  io_out_0_ar_bits_burst,
  output [11:0] io_out_0_ar_bits_user,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [3:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input  [11:0] io_out_0_r_bits_user,
  input         io_out_0_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [63:0] Queue_io_enq_bits_data;
  wire [1:0] Queue_io_enq_bits_resp;
  wire [11:0] Queue_io_enq_bits_user;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [63:0] Queue_io_deq_bits_data;
  wire [1:0] Queue_io_deq_bits_resp;
  wire [11:0] Queue_io_deq_bits_user;
  wire  Queue_io_deq_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [3:0] Queue_1_io_enq_bits_id;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [1:0] Queue_1_io_enq_bits_resp;
  wire [11:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [3:0] Queue_1_io_deq_bits_id;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [1:0] Queue_1_io_deq_bits_resp;
  wire [11:0] Queue_1_io_deq_bits_user;
  wire  Queue_1_io_deq_bits_last;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire [11:0] Queue_2_io_enq_bits_user;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire [11:0] Queue_2_io_deq_bits_user;
  wire  Queue_2_io_deq_bits_last;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [63:0] Queue_3_io_enq_bits_data;
  wire [1:0] Queue_3_io_enq_bits_resp;
  wire [11:0] Queue_3_io_enq_bits_user;
  wire  Queue_3_io_enq_bits_last;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [63:0] Queue_3_io_deq_bits_data;
  wire [1:0] Queue_3_io_deq_bits_resp;
  wire [11:0] Queue_3_io_deq_bits_user;
  wire  Queue_3_io_deq_bits_last;
  reg  _T_380;
  reg [31:0] _RAND_0;
  reg [3:0] _T_382;
  reg [31:0] _RAND_1;
  wire [15:0] _T_385;
  wire [15:0] _T_389;
  reg [3:0] _T_393;
  reg [31:0] _RAND_2;
  wire  _T_395;
  wire  _T_396;
  wire  _T_397;
  wire  _T_398;
  wire  _T_399;
  wire  _T_400;
  wire  _T_401;
  wire  _T_402;
  wire [3:0] _GEN_0;
  wire [4:0] _T_403;
  wire [3:0] _T_404;
  wire [3:0] _GEN_1;
  wire [4:0] _T_405;
  wire [4:0] _T_406;
  wire [3:0] _T_407;
  wire  _T_409;
  wire  _T_411;
  wire  _T_412;
  wire  _T_413;
  wire  _T_415;
  wire  _T_417;
  wire  _T_419;
  wire  _T_420;
  wire  _T_421;
  wire  _T_423;
  wire  _T_425;
  reg [3:0] _T_428;
  reg [31:0] _RAND_3;
  wire  _T_430;
  wire  _T_432;
  wire  _T_433;
  wire  _T_434;
  wire  _T_436;
  wire  _T_437;
  wire [3:0] _GEN_2;
  wire [4:0] _T_438;
  wire [3:0] _T_439;
  wire [3:0] _GEN_3;
  wire [4:0] _T_440;
  wire [4:0] _T_441;
  wire [3:0] _T_442;
  wire  _T_444;
  wire  _T_446;
  wire  _T_447;
  wire  _T_448;
  wire  _T_450;
  wire  _T_452;
  wire  _T_454;
  wire  _T_455;
  wire  _T_456;
  wire  _T_458;
  wire  _T_460;
  reg [3:0] _T_463;
  reg [31:0] _RAND_4;
  wire  _T_465;
  wire  _T_467;
  wire  _T_468;
  wire  _T_469;
  wire  _T_471;
  wire  _T_472;
  wire [3:0] _GEN_4;
  wire [4:0] _T_473;
  wire [3:0] _T_474;
  wire [3:0] _GEN_98;
  wire [4:0] _T_475;
  wire [4:0] _T_476;
  wire [3:0] _T_477;
  wire  _T_479;
  wire  _T_481;
  wire  _T_482;
  wire  _T_483;
  wire  _T_485;
  wire  _T_487;
  wire  _T_489;
  wire  _T_490;
  wire  _T_491;
  wire  _T_493;
  wire  _T_495;
  reg [3:0] _T_498;
  reg [31:0] _RAND_5;
  wire  _T_500;
  wire  _T_502;
  wire  _T_503;
  wire  _T_504;
  wire  _T_506;
  wire  _T_507;
  wire [3:0] _GEN_99;
  wire [4:0] _T_508;
  wire [3:0] _T_509;
  wire [3:0] _GEN_100;
  wire [4:0] _T_510;
  wire [4:0] _T_511;
  wire [3:0] _T_512;
  wire  _T_514;
  wire  _T_516;
  wire  _T_517;
  wire  _T_518;
  wire  _T_520;
  wire  _T_522;
  wire  _T_524;
  wire  _T_525;
  wire  _T_526;
  wire  _T_528;
  wire  _T_530;
  wire [1:0] _T_543;
  wire [1:0] _T_544;
  wire [3:0] _T_545;
  wire [7:0] _T_549;
  wire [15:0] _T_557;
  wire [16:0] _GEN_101;
  wire [16:0] _T_558;
  wire [15:0] _T_559;
  wire [15:0] _T_560;
  wire [17:0] _GEN_102;
  wire [17:0] _T_561;
  wire [15:0] _T_562;
  wire [15:0] _T_563;
  wire [19:0] _GEN_103;
  wire [19:0] _T_564;
  wire [15:0] _T_565;
  wire [15:0] _T_566;
  wire [23:0] _GEN_104;
  wire [23:0] _T_567;
  wire [15:0] _T_568;
  wire [15:0] _T_569;
  wire [16:0] _GEN_105;
  wire [16:0] _T_571;
  wire [16:0] _T_572;
  wire [16:0] _T_573;
  wire  _T_575;
  wire  _T_577;
  wire  _T_578;
  wire  _T_580;
  wire  _T_581;
  wire [15:0] _T_582;
  wire [15:0] _GEN_107;
  wire [15:0] _T_585;
  wire [7:0] _T_586;
  wire [7:0] _T_587;
  wire  _T_589;
  wire [7:0] _T_590;
  wire [3:0] _T_591;
  wire [3:0] _T_592;
  wire  _T_594;
  wire [3:0] _T_595;
  wire [1:0] _T_596;
  wire [1:0] _T_597;
  wire  _T_599;
  wire [1:0] _T_600;
  wire  _T_601;
  wire [1:0] _T_602;
  wire [2:0] _T_603;
  wire [3:0] _T_604;
  wire [4:0] _T_605;
  wire  _GEN_6;
  wire [4:0] _GEN_7;
  wire [3:0] _T_608_0_id;
  wire [63:0] _T_608_0_data;
  wire [1:0] _T_608_0_resp;
  wire [11:0] _T_608_0_user;
  wire  _T_608_0_last;
  wire [3:0] _T_608_1_id;
  wire [63:0] _T_608_1_data;
  wire [1:0] _T_608_1_resp;
  wire [11:0] _T_608_1_user;
  wire  _T_608_1_last;
  wire [3:0] _T_608_2_id;
  wire [63:0] _T_608_2_data;
  wire [1:0] _T_608_2_resp;
  wire [11:0] _T_608_2_user;
  wire  _T_608_2_last;
  wire [3:0] _T_608_3_id;
  wire [63:0] _T_608_3_data;
  wire [1:0] _T_608_3_resp;
  wire [11:0] _T_608_3_user;
  wire  _T_608_3_last;
  wire [3:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [1:0] _GEN_10;
  wire [11:0] _GEN_11;
  wire  _GEN_12;
  wire [3:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [11:0] _GEN_16;
  wire  _GEN_17;
  wire [3:0] _GEN_18;
  wire [63:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [11:0] _GEN_21;
  wire  _GEN_22;
  wire [3:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [1:0] _GEN_25;
  wire [11:0] _GEN_26;
  wire  _GEN_27;
  wire [3:0] _GEN_28;
  wire [63:0] _GEN_29;
  wire [1:0] _GEN_30;
  wire [11:0] _GEN_31;
  wire  _GEN_32;
  wire [3:0] _GEN_33;
  wire [63:0] _GEN_34;
  wire [1:0] _GEN_35;
  wire [11:0] _GEN_36;
  wire  _GEN_37;
  wire [3:0] _GEN_38;
  wire [63:0] _GEN_39;
  wire [1:0] _GEN_40;
  wire [11:0] _GEN_41;
  wire  _GEN_42;
  wire [3:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire [1:0] _GEN_45;
  wire [11:0] _GEN_46;
  wire  _GEN_47;
  wire [3:0] _GEN_48;
  wire [63:0] _GEN_49;
  wire [1:0] _GEN_50;
  wire [11:0] _GEN_51;
  wire  _GEN_52;
  wire [3:0] _GEN_53;
  wire [63:0] _GEN_54;
  wire [1:0] _GEN_55;
  wire [11:0] _GEN_56;
  wire  _GEN_57;
  wire [3:0] _GEN_58;
  wire [63:0] _GEN_59;
  wire [1:0] _GEN_60;
  wire [11:0] _GEN_61;
  wire  _GEN_62;
  wire [3:0] _GEN_63;
  wire [63:0] _GEN_64;
  wire [1:0] _GEN_65;
  wire [11:0] _GEN_66;
  wire  _GEN_67;
  wire [3:0] _GEN_68;
  wire [63:0] _GEN_69;
  wire [1:0] _GEN_70;
  wire [11:0] _GEN_71;
  wire  _GEN_72;
  wire [3:0] _GEN_73;
  wire [63:0] _GEN_74;
  wire [1:0] _GEN_75;
  wire [11:0] _GEN_76;
  wire  _GEN_77;
  wire [3:0] _GEN_78;
  wire [63:0] _GEN_79;
  wire [1:0] _GEN_80;
  wire [11:0] _GEN_81;
  wire  _GEN_82;
  wire  _T_678_0;
  wire  _T_678_1;
  wire  _T_678_2;
  wire  _T_678_3;
  wire  _GEN_83;
  wire  _GEN_84;
  wire  _GEN_85;
  wire  _GEN_86;
  wire  _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire  _GEN_91;
  wire  _GEN_92;
  wire  _GEN_93;
  wire  _GEN_94;
  wire  _GEN_95;
  wire  _GEN_96;
  wire  _GEN_97;
  wire  _T_714;
  wire  _T_715;
  wire  _T_716;
  wire  _T_717;
  Queue_13 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_enq_bits_resp(Queue_io_enq_bits_resp),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_data(Queue_io_deq_bits_data),
    .io_deq_bits_resp(Queue_io_deq_bits_resp),
    .io_deq_bits_user(Queue_io_deq_bits_user),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_13 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_resp(Queue_1_io_enq_bits_resp),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_resp(Queue_1_io_deq_bits_resp),
    .io_deq_bits_user(Queue_1_io_deq_bits_user),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_13 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_enq_bits_user(Queue_2_io_enq_bits_user),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp),
    .io_deq_bits_user(Queue_2_io_deq_bits_user),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  Queue_13 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_data(Queue_3_io_enq_bits_data),
    .io_enq_bits_resp(Queue_3_io_enq_bits_resp),
    .io_enq_bits_user(Queue_3_io_enq_bits_user),
    .io_enq_bits_last(Queue_3_io_enq_bits_last),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_data(Queue_3_io_deq_bits_data),
    .io_deq_bits_resp(Queue_3_io_deq_bits_resp),
    .io_deq_bits_user(Queue_3_io_deq_bits_user),
    .io_deq_bits_last(Queue_3_io_deq_bits_last)
  );
  assign io_in_0_aw_ready = io_out_0_aw_ready;
  assign io_in_0_w_ready = io_out_0_w_ready;
  assign io_in_0_b_valid = io_out_0_b_valid;
  assign io_in_0_b_bits_id = io_out_0_b_bits_id;
  assign io_in_0_b_bits_resp = io_out_0_b_bits_resp;
  assign io_in_0_b_bits_user = io_out_0_b_bits_user;
  assign io_in_0_ar_ready = io_out_0_ar_ready;
  assign io_in_0_r_valid = _T_380;
  assign io_in_0_r_bits_id = _GEN_78;
  assign io_in_0_r_bits_data = _GEN_79;
  assign io_in_0_r_bits_resp = _GEN_80;
  assign io_in_0_r_bits_user = _GEN_81;
  assign io_in_0_r_bits_last = _GEN_82;
  assign io_out_0_aw_valid = io_in_0_aw_valid;
  assign io_out_0_aw_bits_id = io_in_0_aw_bits_id;
  assign io_out_0_aw_bits_addr = io_in_0_aw_bits_addr;
  assign io_out_0_aw_bits_len = io_in_0_aw_bits_len;
  assign io_out_0_aw_bits_size = io_in_0_aw_bits_size;
  assign io_out_0_aw_bits_burst = io_in_0_aw_bits_burst;
  assign io_out_0_aw_bits_user = io_in_0_aw_bits_user;
  assign io_out_0_w_valid = io_in_0_w_valid;
  assign io_out_0_w_bits_data = io_in_0_w_bits_data;
  assign io_out_0_w_bits_strb = io_in_0_w_bits_strb;
  assign io_out_0_w_bits_last = io_in_0_w_bits_last;
  assign io_out_0_b_ready = io_in_0_b_ready;
  assign io_out_0_ar_valid = io_in_0_ar_valid;
  assign io_out_0_ar_bits_id = io_in_0_ar_bits_id;
  assign io_out_0_ar_bits_addr = io_in_0_ar_bits_addr;
  assign io_out_0_ar_bits_len = io_in_0_ar_bits_len;
  assign io_out_0_ar_bits_size = io_in_0_ar_bits_size;
  assign io_out_0_ar_bits_burst = io_in_0_ar_bits_burst;
  assign io_out_0_ar_bits_user = io_in_0_ar_bits_user;
  assign io_out_0_r_ready = _GEN_97;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_714;
  assign Queue_io_enq_bits_id = io_out_0_r_bits_id;
  assign Queue_io_enq_bits_data = io_out_0_r_bits_data;
  assign Queue_io_enq_bits_resp = io_out_0_r_bits_resp;
  assign Queue_io_enq_bits_user = io_out_0_r_bits_user;
  assign Queue_io_enq_bits_last = io_out_0_r_bits_last;
  assign Queue_io_deq_ready = _T_401;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_715;
  assign Queue_1_io_enq_bits_id = io_out_0_r_bits_id;
  assign Queue_1_io_enq_bits_data = io_out_0_r_bits_data;
  assign Queue_1_io_enq_bits_resp = io_out_0_r_bits_resp;
  assign Queue_1_io_enq_bits_user = io_out_0_r_bits_user;
  assign Queue_1_io_enq_bits_last = io_out_0_r_bits_last;
  assign Queue_1_io_deq_ready = _T_436;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = _T_716;
  assign Queue_2_io_enq_bits_id = io_out_0_r_bits_id;
  assign Queue_2_io_enq_bits_data = io_out_0_r_bits_data;
  assign Queue_2_io_enq_bits_resp = io_out_0_r_bits_resp;
  assign Queue_2_io_enq_bits_user = io_out_0_r_bits_user;
  assign Queue_2_io_enq_bits_last = io_out_0_r_bits_last;
  assign Queue_2_io_deq_ready = _T_471;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = _T_717;
  assign Queue_3_io_enq_bits_id = io_out_0_r_bits_id;
  assign Queue_3_io_enq_bits_data = io_out_0_r_bits_data;
  assign Queue_3_io_enq_bits_resp = io_out_0_r_bits_resp;
  assign Queue_3_io_enq_bits_user = io_out_0_r_bits_user;
  assign Queue_3_io_enq_bits_last = io_out_0_r_bits_last;
  assign Queue_3_io_deq_ready = _T_506;
  assign _T_385 = 16'h1 << _T_382;
  assign _T_389 = 16'h1 << io_out_0_r_bits_id;
  assign _T_395 = _T_389[0];
  assign _T_396 = io_out_0_r_ready & io_out_0_r_valid;
  assign _T_397 = _T_395 & _T_396;
  assign _T_398 = _T_397 & io_out_0_r_bits_last;
  assign _T_399 = _T_385[0];
  assign _T_400 = io_in_0_r_ready & io_in_0_r_valid;
  assign _T_401 = _T_399 & _T_400;
  assign _T_402 = _T_401 & io_in_0_r_bits_last;
  assign _GEN_0 = {{3'd0}, _T_398};
  assign _T_403 = _T_393 + _GEN_0;
  assign _T_404 = _T_403[3:0];
  assign _GEN_1 = {{3'd0}, _T_402};
  assign _T_405 = _T_404 - _GEN_1;
  assign _T_406 = $unsigned(_T_405);
  assign _T_407 = _T_406[3:0];
  assign _T_409 = _T_402 == 1'h0;
  assign _T_411 = _T_393 != 4'h0;
  assign _T_412 = _T_409 | _T_411;
  assign _T_413 = _T_412 | reset;
  assign _T_415 = _T_413 == 1'h0;
  assign _T_417 = _T_398 == 1'h0;
  assign _T_419 = _T_393 != 4'h8;
  assign _T_420 = _T_417 | _T_419;
  assign _T_421 = _T_420 | reset;
  assign _T_423 = _T_421 == 1'h0;
  assign _T_425 = _T_407 != 4'h0;
  assign _T_430 = _T_389[1];
  assign _T_432 = _T_430 & _T_396;
  assign _T_433 = _T_432 & io_out_0_r_bits_last;
  assign _T_434 = _T_385[1];
  assign _T_436 = _T_434 & _T_400;
  assign _T_437 = _T_436 & io_in_0_r_bits_last;
  assign _GEN_2 = {{3'd0}, _T_433};
  assign _T_438 = _T_428 + _GEN_2;
  assign _T_439 = _T_438[3:0];
  assign _GEN_3 = {{3'd0}, _T_437};
  assign _T_440 = _T_439 - _GEN_3;
  assign _T_441 = $unsigned(_T_440);
  assign _T_442 = _T_441[3:0];
  assign _T_444 = _T_437 == 1'h0;
  assign _T_446 = _T_428 != 4'h0;
  assign _T_447 = _T_444 | _T_446;
  assign _T_448 = _T_447 | reset;
  assign _T_450 = _T_448 == 1'h0;
  assign _T_452 = _T_433 == 1'h0;
  assign _T_454 = _T_428 != 4'h8;
  assign _T_455 = _T_452 | _T_454;
  assign _T_456 = _T_455 | reset;
  assign _T_458 = _T_456 == 1'h0;
  assign _T_460 = _T_442 != 4'h0;
  assign _T_465 = _T_389[2];
  assign _T_467 = _T_465 & _T_396;
  assign _T_468 = _T_467 & io_out_0_r_bits_last;
  assign _T_469 = _T_385[2];
  assign _T_471 = _T_469 & _T_400;
  assign _T_472 = _T_471 & io_in_0_r_bits_last;
  assign _GEN_4 = {{3'd0}, _T_468};
  assign _T_473 = _T_463 + _GEN_4;
  assign _T_474 = _T_473[3:0];
  assign _GEN_98 = {{3'd0}, _T_472};
  assign _T_475 = _T_474 - _GEN_98;
  assign _T_476 = $unsigned(_T_475);
  assign _T_477 = _T_476[3:0];
  assign _T_479 = _T_472 == 1'h0;
  assign _T_481 = _T_463 != 4'h0;
  assign _T_482 = _T_479 | _T_481;
  assign _T_483 = _T_482 | reset;
  assign _T_485 = _T_483 == 1'h0;
  assign _T_487 = _T_468 == 1'h0;
  assign _T_489 = _T_463 != 4'h8;
  assign _T_490 = _T_487 | _T_489;
  assign _T_491 = _T_490 | reset;
  assign _T_493 = _T_491 == 1'h0;
  assign _T_495 = _T_477 != 4'h0;
  assign _T_500 = _T_389[3];
  assign _T_502 = _T_500 & _T_396;
  assign _T_503 = _T_502 & io_out_0_r_bits_last;
  assign _T_504 = _T_385[3];
  assign _T_506 = _T_504 & _T_400;
  assign _T_507 = _T_506 & io_in_0_r_bits_last;
  assign _GEN_99 = {{3'd0}, _T_503};
  assign _T_508 = _T_498 + _GEN_99;
  assign _T_509 = _T_508[3:0];
  assign _GEN_100 = {{3'd0}, _T_507};
  assign _T_510 = _T_509 - _GEN_100;
  assign _T_511 = $unsigned(_T_510);
  assign _T_512 = _T_511[3:0];
  assign _T_514 = _T_507 == 1'h0;
  assign _T_516 = _T_498 != 4'h0;
  assign _T_517 = _T_514 | _T_516;
  assign _T_518 = _T_517 | reset;
  assign _T_520 = _T_518 == 1'h0;
  assign _T_522 = _T_503 == 1'h0;
  assign _T_524 = _T_498 != 4'h8;
  assign _T_525 = _T_522 | _T_524;
  assign _T_526 = _T_525 | reset;
  assign _T_528 = _T_526 == 1'h0;
  assign _T_530 = _T_512 != 4'h0;
  assign _T_543 = {_T_460,_T_425};
  assign _T_544 = {_T_530,_T_495};
  assign _T_545 = {_T_544,_T_543};
  assign _T_549 = {4'h0,_T_545};
  assign _T_557 = {8'h0,_T_549};
  assign _GEN_101 = {{1'd0}, _T_557};
  assign _T_558 = _GEN_101 << 1;
  assign _T_559 = _T_558[15:0];
  assign _T_560 = _T_557 | _T_559;
  assign _GEN_102 = {{2'd0}, _T_560};
  assign _T_561 = _GEN_102 << 2;
  assign _T_562 = _T_561[15:0];
  assign _T_563 = _T_560 | _T_562;
  assign _GEN_103 = {{4'd0}, _T_563};
  assign _T_564 = _GEN_103 << 4;
  assign _T_565 = _T_564[15:0];
  assign _T_566 = _T_563 | _T_565;
  assign _GEN_104 = {{8'd0}, _T_566};
  assign _T_567 = _GEN_104 << 8;
  assign _T_568 = _T_567[15:0];
  assign _T_569 = _T_566 | _T_568;
  assign _GEN_105 = {{1'd0}, _T_569};
  assign _T_571 = _GEN_105 << 1;
  assign _T_572 = ~ _T_571;
  assign _T_573 = _GEN_101 & _T_572;
  assign _T_575 = _T_380 == 1'h0;
  assign _T_577 = _T_400 & io_in_0_r_bits_last;
  assign _T_578 = _T_575 | _T_577;
  assign _T_580 = _T_557 != 16'h0;
  assign _T_581 = _T_573[16];
  assign _T_582 = _T_573[15:0];
  assign _GEN_107 = {{15'd0}, _T_581};
  assign _T_585 = _GEN_107 | _T_582;
  assign _T_586 = _T_585[15:8];
  assign _T_587 = _T_585[7:0];
  assign _T_589 = _T_586 != 8'h0;
  assign _T_590 = _T_586 | _T_587;
  assign _T_591 = _T_590[7:4];
  assign _T_592 = _T_590[3:0];
  assign _T_594 = _T_591 != 4'h0;
  assign _T_595 = _T_591 | _T_592;
  assign _T_596 = _T_595[3:2];
  assign _T_597 = _T_595[1:0];
  assign _T_599 = _T_596 != 2'h0;
  assign _T_600 = _T_596 | _T_597;
  assign _T_601 = _T_600[1];
  assign _T_602 = {_T_599,_T_601};
  assign _T_603 = {_T_594,_T_602};
  assign _T_604 = {_T_589,_T_603};
  assign _T_605 = {_T_581,_T_604};
  assign _GEN_6 = _T_578 ? _T_580 : _T_380;
  assign _GEN_7 = _T_578 ? _T_605 : {{1'd0}, _T_382};
  assign _T_608_0_id = Queue_io_deq_bits_id;
  assign _T_608_0_data = Queue_io_deq_bits_data;
  assign _T_608_0_resp = Queue_io_deq_bits_resp;
  assign _T_608_0_user = Queue_io_deq_bits_user;
  assign _T_608_0_last = Queue_io_deq_bits_last;
  assign _T_608_1_id = Queue_1_io_deq_bits_id;
  assign _T_608_1_data = Queue_1_io_deq_bits_data;
  assign _T_608_1_resp = Queue_1_io_deq_bits_resp;
  assign _T_608_1_user = Queue_1_io_deq_bits_user;
  assign _T_608_1_last = Queue_1_io_deq_bits_last;
  assign _T_608_2_id = Queue_2_io_deq_bits_id;
  assign _T_608_2_data = Queue_2_io_deq_bits_data;
  assign _T_608_2_resp = Queue_2_io_deq_bits_resp;
  assign _T_608_2_user = Queue_2_io_deq_bits_user;
  assign _T_608_2_last = Queue_2_io_deq_bits_last;
  assign _T_608_3_id = Queue_3_io_deq_bits_id;
  assign _T_608_3_data = Queue_3_io_deq_bits_data;
  assign _T_608_3_resp = Queue_3_io_deq_bits_resp;
  assign _T_608_3_user = Queue_3_io_deq_bits_user;
  assign _T_608_3_last = Queue_3_io_deq_bits_last;
  assign _GEN_8 = 4'h1 == _T_382 ? _T_608_1_id : _T_608_0_id;
  assign _GEN_9 = 4'h1 == _T_382 ? _T_608_1_data : _T_608_0_data;
  assign _GEN_10 = 4'h1 == _T_382 ? _T_608_1_resp : _T_608_0_resp;
  assign _GEN_11 = 4'h1 == _T_382 ? _T_608_1_user : _T_608_0_user;
  assign _GEN_12 = 4'h1 == _T_382 ? _T_608_1_last : _T_608_0_last;
  assign _GEN_13 = 4'h2 == _T_382 ? _T_608_2_id : _GEN_8;
  assign _GEN_14 = 4'h2 == _T_382 ? _T_608_2_data : _GEN_9;
  assign _GEN_15 = 4'h2 == _T_382 ? _T_608_2_resp : _GEN_10;
  assign _GEN_16 = 4'h2 == _T_382 ? _T_608_2_user : _GEN_11;
  assign _GEN_17 = 4'h2 == _T_382 ? _T_608_2_last : _GEN_12;
  assign _GEN_18 = 4'h3 == _T_382 ? _T_608_3_id : _GEN_13;
  assign _GEN_19 = 4'h3 == _T_382 ? _T_608_3_data : _GEN_14;
  assign _GEN_20 = 4'h3 == _T_382 ? _T_608_3_resp : _GEN_15;
  assign _GEN_21 = 4'h3 == _T_382 ? _T_608_3_user : _GEN_16;
  assign _GEN_22 = 4'h3 == _T_382 ? _T_608_3_last : _GEN_17;
  assign _GEN_23 = 4'h4 == _T_382 ? 4'h0 : _GEN_18;
  assign _GEN_24 = 4'h4 == _T_382 ? 64'h0 : _GEN_19;
  assign _GEN_25 = 4'h4 == _T_382 ? 2'h0 : _GEN_20;
  assign _GEN_26 = 4'h4 == _T_382 ? 12'h0 : _GEN_21;
  assign _GEN_27 = 4'h4 == _T_382 ? 1'h0 : _GEN_22;
  assign _GEN_28 = 4'h5 == _T_382 ? 4'h0 : _GEN_23;
  assign _GEN_29 = 4'h5 == _T_382 ? 64'h0 : _GEN_24;
  assign _GEN_30 = 4'h5 == _T_382 ? 2'h0 : _GEN_25;
  assign _GEN_31 = 4'h5 == _T_382 ? 12'h0 : _GEN_26;
  assign _GEN_32 = 4'h5 == _T_382 ? 1'h0 : _GEN_27;
  assign _GEN_33 = 4'h6 == _T_382 ? 4'h0 : _GEN_28;
  assign _GEN_34 = 4'h6 == _T_382 ? 64'h0 : _GEN_29;
  assign _GEN_35 = 4'h6 == _T_382 ? 2'h0 : _GEN_30;
  assign _GEN_36 = 4'h6 == _T_382 ? 12'h0 : _GEN_31;
  assign _GEN_37 = 4'h6 == _T_382 ? 1'h0 : _GEN_32;
  assign _GEN_38 = 4'h7 == _T_382 ? 4'h0 : _GEN_33;
  assign _GEN_39 = 4'h7 == _T_382 ? 64'h0 : _GEN_34;
  assign _GEN_40 = 4'h7 == _T_382 ? 2'h0 : _GEN_35;
  assign _GEN_41 = 4'h7 == _T_382 ? 12'h0 : _GEN_36;
  assign _GEN_42 = 4'h7 == _T_382 ? 1'h0 : _GEN_37;
  assign _GEN_43 = 4'h8 == _T_382 ? 4'h0 : _GEN_38;
  assign _GEN_44 = 4'h8 == _T_382 ? 64'h0 : _GEN_39;
  assign _GEN_45 = 4'h8 == _T_382 ? 2'h0 : _GEN_40;
  assign _GEN_46 = 4'h8 == _T_382 ? 12'h0 : _GEN_41;
  assign _GEN_47 = 4'h8 == _T_382 ? 1'h0 : _GEN_42;
  assign _GEN_48 = 4'h9 == _T_382 ? 4'h0 : _GEN_43;
  assign _GEN_49 = 4'h9 == _T_382 ? 64'h0 : _GEN_44;
  assign _GEN_50 = 4'h9 == _T_382 ? 2'h0 : _GEN_45;
  assign _GEN_51 = 4'h9 == _T_382 ? 12'h0 : _GEN_46;
  assign _GEN_52 = 4'h9 == _T_382 ? 1'h0 : _GEN_47;
  assign _GEN_53 = 4'ha == _T_382 ? 4'h0 : _GEN_48;
  assign _GEN_54 = 4'ha == _T_382 ? 64'h0 : _GEN_49;
  assign _GEN_55 = 4'ha == _T_382 ? 2'h0 : _GEN_50;
  assign _GEN_56 = 4'ha == _T_382 ? 12'h0 : _GEN_51;
  assign _GEN_57 = 4'ha == _T_382 ? 1'h0 : _GEN_52;
  assign _GEN_58 = 4'hb == _T_382 ? 4'h0 : _GEN_53;
  assign _GEN_59 = 4'hb == _T_382 ? 64'h0 : _GEN_54;
  assign _GEN_60 = 4'hb == _T_382 ? 2'h0 : _GEN_55;
  assign _GEN_61 = 4'hb == _T_382 ? 12'h0 : _GEN_56;
  assign _GEN_62 = 4'hb == _T_382 ? 1'h0 : _GEN_57;
  assign _GEN_63 = 4'hc == _T_382 ? 4'h0 : _GEN_58;
  assign _GEN_64 = 4'hc == _T_382 ? 64'h0 : _GEN_59;
  assign _GEN_65 = 4'hc == _T_382 ? 2'h0 : _GEN_60;
  assign _GEN_66 = 4'hc == _T_382 ? 12'h0 : _GEN_61;
  assign _GEN_67 = 4'hc == _T_382 ? 1'h0 : _GEN_62;
  assign _GEN_68 = 4'hd == _T_382 ? 4'h0 : _GEN_63;
  assign _GEN_69 = 4'hd == _T_382 ? 64'h0 : _GEN_64;
  assign _GEN_70 = 4'hd == _T_382 ? 2'h0 : _GEN_65;
  assign _GEN_71 = 4'hd == _T_382 ? 12'h0 : _GEN_66;
  assign _GEN_72 = 4'hd == _T_382 ? 1'h0 : _GEN_67;
  assign _GEN_73 = 4'he == _T_382 ? 4'h0 : _GEN_68;
  assign _GEN_74 = 4'he == _T_382 ? 64'h0 : _GEN_69;
  assign _GEN_75 = 4'he == _T_382 ? 2'h0 : _GEN_70;
  assign _GEN_76 = 4'he == _T_382 ? 12'h0 : _GEN_71;
  assign _GEN_77 = 4'he == _T_382 ? 1'h0 : _GEN_72;
  assign _GEN_78 = 4'hf == _T_382 ? 4'h0 : _GEN_73;
  assign _GEN_79 = 4'hf == _T_382 ? 64'h0 : _GEN_74;
  assign _GEN_80 = 4'hf == _T_382 ? 2'h0 : _GEN_75;
  assign _GEN_81 = 4'hf == _T_382 ? 12'h0 : _GEN_76;
  assign _GEN_82 = 4'hf == _T_382 ? 1'h0 : _GEN_77;
  assign _T_678_0 = Queue_io_enq_ready;
  assign _T_678_1 = Queue_1_io_enq_ready;
  assign _T_678_2 = Queue_2_io_enq_ready;
  assign _T_678_3 = Queue_3_io_enq_ready;
  assign _GEN_83 = 4'h1 == io_out_0_r_bits_id ? _T_678_1 : _T_678_0;
  assign _GEN_84 = 4'h2 == io_out_0_r_bits_id ? _T_678_2 : _GEN_83;
  assign _GEN_85 = 4'h3 == io_out_0_r_bits_id ? _T_678_3 : _GEN_84;
  assign _GEN_86 = 4'h4 == io_out_0_r_bits_id ? 1'h0 : _GEN_85;
  assign _GEN_87 = 4'h5 == io_out_0_r_bits_id ? 1'h0 : _GEN_86;
  assign _GEN_88 = 4'h6 == io_out_0_r_bits_id ? 1'h0 : _GEN_87;
  assign _GEN_89 = 4'h7 == io_out_0_r_bits_id ? 1'h0 : _GEN_88;
  assign _GEN_90 = 4'h8 == io_out_0_r_bits_id ? 1'h0 : _GEN_89;
  assign _GEN_91 = 4'h9 == io_out_0_r_bits_id ? 1'h0 : _GEN_90;
  assign _GEN_92 = 4'ha == io_out_0_r_bits_id ? 1'h0 : _GEN_91;
  assign _GEN_93 = 4'hb == io_out_0_r_bits_id ? 1'h0 : _GEN_92;
  assign _GEN_94 = 4'hc == io_out_0_r_bits_id ? 1'h0 : _GEN_93;
  assign _GEN_95 = 4'hd == io_out_0_r_bits_id ? 1'h0 : _GEN_94;
  assign _GEN_96 = 4'he == io_out_0_r_bits_id ? 1'h0 : _GEN_95;
  assign _GEN_97 = 4'hf == io_out_0_r_bits_id ? 1'h0 : _GEN_96;
  assign _T_714 = _T_395 & io_out_0_r_valid;
  assign _T_715 = _T_430 & io_out_0_r_valid;
  assign _T_716 = _T_465 & io_out_0_r_valid;
  assign _T_717 = _T_500 & io_out_0_r_valid;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_380 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_382 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_393 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_428 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_463 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_498 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_380 <= 1'h0;
    end else begin
      if (_T_578) begin
        _T_380 <= _T_580;
      end
    end
    _T_382 <= _GEN_7[3:0];
    if (reset) begin
      _T_393 <= 4'h0;
    end else begin
      _T_393 <= _T_407;
    end
    if (reset) begin
      _T_428 <= 4'h0;
    end else begin
      _T_428 <= _T_442;
    end
    if (reset) begin
      _T_463 <= 4'h0;
    end else begin
      _T_463 <= _T_477;
    end
    if (reset) begin
      _T_498 <= 4'h0;
    end else begin
      _T_498 <= _T_512;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_415) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:75 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_415) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_423) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:76 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_423) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_450) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:75 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_450) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_458) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:76 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_458) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_485) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:75 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_485) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_493) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:76 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_493) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_520) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:75 assert (!dec || count =/= UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_520) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_528) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Deinterleaver.scala:76 assert (!inc || count =/= UInt(beats))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_528) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_17(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [11:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [11:0] io_deq_bits
);
  reg [11:0] ram [0:0];
  reg [31:0] _RAND_0;
  wire [11:0] ram__T_35_data;
  wire  ram__T_35_addr;
  wire [11:0] ram__T_26_data;
  wire  ram__T_26_addr;
  wire  ram__T_26_mask;
  wire  ram__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_1;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_4;
  wire  _T_31;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _T_31;
  assign io_deq_bits = ram__T_35_data;
  assign ram__T_35_addr = 1'h0;
  assign ram__T_35_data = ram[ram__T_35_addr];
  assign ram__T_26_data = io_enq_bits;
  assign ram__T_26_addr = 1'h0;
  assign ram__T_26_mask = _T_21;
  assign ram__T_26_en = _T_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _T_21 != _T_23;
  assign _GEN_4 = _T_29 ? _T_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  maybe_full = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_26_en & ram__T_26_mask) begin
      ram[ram__T_26_addr] <= ram__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        maybe_full <= _T_21;
      end
    end
  end
endmodule
module Queue_19(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [11:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [11:0] io_deq_bits
);
  reg [11:0] ram [0:7];
  reg [31:0] _RAND_0;
  wire [11:0] ram__T_43_data;
  wire [2:0] ram__T_43_addr;
  wire [11:0] ram__T_29_data;
  wire [2:0] ram__T_29_addr;
  wire  ram__T_29_mask;
  wire  ram__T_29_en;
  reg [2:0] value;
  reg [31:0] _RAND_1;
  reg [2:0] value_1;
  reg [31:0] _RAND_2;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [3:0] _T_32;
  wire [2:0] _T_33;
  wire [2:0] _GEN_4;
  wire [3:0] _T_36;
  wire [2:0] _T_37;
  wire [2:0] _GEN_5;
  wire  _T_38;
  wire  _GEN_6;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits = ram__T_43_data;
  assign ram__T_43_addr = value_1;
  assign ram__T_43_data = ram[ram__T_43_addr];
  assign ram__T_29_data = io_enq_bits;
  assign ram__T_29_addr = value;
  assign ram__T_29_mask = _T_25;
  assign ram__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 3'h1;
  assign _T_33 = _T_32[2:0];
  assign _GEN_4 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 3'h1;
  assign _T_37 = _T_36[2:0];
  assign _GEN_5 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_6 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ram[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  value = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value_1 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_29_en & ram__T_29_mask) begin
      ram[ram__T_29_addr] <= ram__T_29_data;
    end
    if (reset) begin
      value <= 3'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module AXI4UserYanker(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [3:0]  io_in_0_aw_bits_id,
  input  [30:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  input  [11:0] io_in_0_aw_bits_user,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [3:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output [11:0] io_in_0_b_bits_user,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [3:0]  io_in_0_ar_bits_id,
  input  [30:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input  [11:0] io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [3:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output [11:0] io_in_0_r_bits_user,
  output        io_in_0_r_bits_last,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [3:0]  io_out_0_aw_bits_id,
  output [30:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [1:0]  io_out_0_aw_bits_burst,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [3:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [3:0]  io_out_0_ar_bits_id,
  output [30:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [1:0]  io_out_0_ar_bits_burst,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [3:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input         io_out_0_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [11:0] Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [11:0] Queue_io_deq_bits;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [11:0] Queue_1_io_enq_bits;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [11:0] Queue_1_io_deq_bits;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [11:0] Queue_2_io_enq_bits;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [11:0] Queue_2_io_deq_bits;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [11:0] Queue_3_io_enq_bits;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [11:0] Queue_3_io_deq_bits;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [11:0] Queue_4_io_enq_bits;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [11:0] Queue_4_io_deq_bits;
  wire  Queue_5_clock;
  wire  Queue_5_reset;
  wire  Queue_5_io_enq_ready;
  wire  Queue_5_io_enq_valid;
  wire [11:0] Queue_5_io_enq_bits;
  wire  Queue_5_io_deq_ready;
  wire  Queue_5_io_deq_valid;
  wire [11:0] Queue_5_io_deq_bits;
  wire  Queue_6_clock;
  wire  Queue_6_reset;
  wire  Queue_6_io_enq_ready;
  wire  Queue_6_io_enq_valid;
  wire [11:0] Queue_6_io_enq_bits;
  wire  Queue_6_io_deq_ready;
  wire  Queue_6_io_deq_valid;
  wire [11:0] Queue_6_io_deq_bits;
  wire  Queue_7_clock;
  wire  Queue_7_reset;
  wire  Queue_7_io_enq_ready;
  wire  Queue_7_io_enq_valid;
  wire [11:0] Queue_7_io_enq_bits;
  wire  Queue_7_io_deq_ready;
  wire  Queue_7_io_deq_valid;
  wire [11:0] Queue_7_io_deq_bits;
  wire  _T_700_0;
  wire  _T_700_1;
  wire  _T_700_2;
  wire  _T_700_3;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire  _GEN_20;
  wire  _GEN_21;
  wire  _GEN_22;
  wire  _T_720;
  wire  _T_721;
  wire  _T_724_0;
  wire  _T_724_1;
  wire  _T_724_2;
  wire  _T_724_3;
  wire [11:0] _T_746_0;
  wire [11:0] _T_746_1;
  wire [11:0] _T_746_2;
  wire [11:0] _T_746_3;
  wire  _T_767;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire  _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire  _GEN_35;
  wire  _GEN_36;
  wire  _GEN_37;
  wire  _T_768;
  wire  _T_769;
  wire  _T_771;
  wire [11:0] _GEN_38;
  wire [11:0] _GEN_39;
  wire [11:0] _GEN_40;
  wire [11:0] _GEN_41;
  wire [11:0] _GEN_42;
  wire [11:0] _GEN_43;
  wire [11:0] _GEN_44;
  wire [11:0] _GEN_45;
  wire [11:0] _GEN_46;
  wire [11:0] _GEN_47;
  wire [11:0] _GEN_48;
  wire [11:0] _GEN_49;
  wire [11:0] _GEN_50;
  wire [11:0] _GEN_51;
  wire [11:0] _GEN_52;
  wire [15:0] _T_774;
  wire  _T_776;
  wire  _T_777;
  wire  _T_778;
  wire  _T_779;
  wire [15:0] _T_794;
  wire  _T_796;
  wire  _T_797;
  wire  _T_798;
  wire  _T_799;
  wire  _T_812;
  wire  _T_813;
  wire  _T_814;
  wire  _T_815;
  wire  _T_816;
  wire  _T_818;
  wire  _T_819;
  wire  _T_821;
  wire  _T_823;
  wire  _T_824;
  wire  _T_826;
  wire  _T_828;
  wire  _T_829;
  wire  _T_831;
  wire  _T_894_0;
  wire  _T_894_1;
  wire  _T_894_2;
  wire  _T_894_3;
  wire  _GEN_53;
  wire  _GEN_54;
  wire  _GEN_55;
  wire  _GEN_56;
  wire  _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire  _GEN_60;
  wire  _GEN_61;
  wire  _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire  _GEN_65;
  wire  _GEN_66;
  wire  _GEN_67;
  wire  _T_914;
  wire  _T_915;
  wire  _T_918_0;
  wire  _T_918_1;
  wire  _T_918_2;
  wire  _T_918_3;
  wire [11:0] _T_940_0;
  wire [11:0] _T_940_1;
  wire [11:0] _T_940_2;
  wire [11:0] _T_940_3;
  wire  _T_961;
  wire  _GEN_68;
  wire  _GEN_69;
  wire  _GEN_70;
  wire  _GEN_71;
  wire  _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire  _GEN_75;
  wire  _GEN_76;
  wire  _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire  _T_962;
  wire  _T_963;
  wire  _T_965;
  wire [11:0] _GEN_83;
  wire [11:0] _GEN_84;
  wire [11:0] _GEN_85;
  wire [11:0] _GEN_86;
  wire [11:0] _GEN_87;
  wire [11:0] _GEN_88;
  wire [11:0] _GEN_89;
  wire [11:0] _GEN_90;
  wire [11:0] _GEN_91;
  wire [11:0] _GEN_92;
  wire [11:0] _GEN_93;
  wire [11:0] _GEN_94;
  wire [11:0] _GEN_95;
  wire [11:0] _GEN_96;
  wire [11:0] _GEN_97;
  wire [15:0] _T_968;
  wire  _T_970;
  wire  _T_971;
  wire  _T_972;
  wire  _T_973;
  wire [15:0] _T_988;
  wire  _T_990;
  wire  _T_991;
  wire  _T_992;
  wire  _T_993;
  wire  _T_1006;
  wire  _T_1007;
  wire  _T_1008;
  wire  _T_1009;
  wire  _T_1011;
  wire  _T_1013;
  wire  _T_1015;
  wire  _T_1017;
  wire  _T_1019;
  wire  _T_1021;
  Queue_17 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_17 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_19 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_19 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  Queue_17 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits(Queue_4_io_enq_bits),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits(Queue_4_io_deq_bits)
  );
  Queue_17 Queue_5 (
    .clock(Queue_5_clock),
    .reset(Queue_5_reset),
    .io_enq_ready(Queue_5_io_enq_ready),
    .io_enq_valid(Queue_5_io_enq_valid),
    .io_enq_bits(Queue_5_io_enq_bits),
    .io_deq_ready(Queue_5_io_deq_ready),
    .io_deq_valid(Queue_5_io_deq_valid),
    .io_deq_bits(Queue_5_io_deq_bits)
  );
  Queue_19 Queue_6 (
    .clock(Queue_6_clock),
    .reset(Queue_6_reset),
    .io_enq_ready(Queue_6_io_enq_ready),
    .io_enq_valid(Queue_6_io_enq_valid),
    .io_enq_bits(Queue_6_io_enq_bits),
    .io_deq_ready(Queue_6_io_deq_ready),
    .io_deq_valid(Queue_6_io_deq_valid),
    .io_deq_bits(Queue_6_io_deq_bits)
  );
  Queue_19 Queue_7 (
    .clock(Queue_7_clock),
    .reset(Queue_7_reset),
    .io_enq_ready(Queue_7_io_enq_ready),
    .io_enq_valid(Queue_7_io_enq_valid),
    .io_enq_bits(Queue_7_io_enq_bits),
    .io_deq_ready(Queue_7_io_deq_ready),
    .io_deq_valid(Queue_7_io_deq_valid),
    .io_deq_bits(Queue_7_io_deq_bits)
  );
  assign io_in_0_aw_ready = _T_914;
  assign io_in_0_w_ready = io_out_0_w_ready;
  assign io_in_0_b_valid = io_out_0_b_valid;
  assign io_in_0_b_bits_id = io_out_0_b_bits_id;
  assign io_in_0_b_bits_resp = io_out_0_b_bits_resp;
  assign io_in_0_b_bits_user = _GEN_97;
  assign io_in_0_ar_ready = _T_720;
  assign io_in_0_r_valid = io_out_0_r_valid;
  assign io_in_0_r_bits_id = io_out_0_r_bits_id;
  assign io_in_0_r_bits_data = io_out_0_r_bits_data;
  assign io_in_0_r_bits_resp = io_out_0_r_bits_resp;
  assign io_in_0_r_bits_user = _GEN_52;
  assign io_in_0_r_bits_last = io_out_0_r_bits_last;
  assign io_out_0_aw_valid = _T_915;
  assign io_out_0_aw_bits_id = io_in_0_aw_bits_id;
  assign io_out_0_aw_bits_addr = io_in_0_aw_bits_addr;
  assign io_out_0_aw_bits_len = io_in_0_aw_bits_len;
  assign io_out_0_aw_bits_size = io_in_0_aw_bits_size;
  assign io_out_0_aw_bits_burst = io_in_0_aw_bits_burst;
  assign io_out_0_w_valid = io_in_0_w_valid;
  assign io_out_0_w_bits_data = io_in_0_w_bits_data;
  assign io_out_0_w_bits_strb = io_in_0_w_bits_strb;
  assign io_out_0_w_bits_last = io_in_0_w_bits_last;
  assign io_out_0_b_ready = io_in_0_b_ready;
  assign io_out_0_ar_valid = _T_721;
  assign io_out_0_ar_bits_id = io_in_0_ar_bits_id;
  assign io_out_0_ar_bits_addr = io_in_0_ar_bits_addr;
  assign io_out_0_ar_bits_len = io_in_0_ar_bits_len;
  assign io_out_0_ar_bits_size = io_in_0_ar_bits_size;
  assign io_out_0_ar_bits_burst = io_in_0_ar_bits_burst;
  assign io_out_0_r_ready = io_in_0_r_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_816;
  assign Queue_io_enq_bits = io_in_0_ar_bits_user;
  assign Queue_io_deq_ready = _T_814;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_821;
  assign Queue_1_io_enq_bits = io_in_0_ar_bits_user;
  assign Queue_1_io_deq_ready = _T_819;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = _T_826;
  assign Queue_2_io_enq_bits = io_in_0_ar_bits_user;
  assign Queue_2_io_deq_ready = _T_824;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = _T_831;
  assign Queue_3_io_enq_bits = io_in_0_ar_bits_user;
  assign Queue_3_io_deq_ready = _T_829;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = _T_1009;
  assign Queue_4_io_enq_bits = io_in_0_aw_bits_user;
  assign Queue_4_io_deq_ready = _T_1007;
  assign Queue_5_clock = clock;
  assign Queue_5_reset = reset;
  assign Queue_5_io_enq_valid = _T_1013;
  assign Queue_5_io_enq_bits = io_in_0_aw_bits_user;
  assign Queue_5_io_deq_ready = _T_1011;
  assign Queue_6_clock = clock;
  assign Queue_6_reset = reset;
  assign Queue_6_io_enq_valid = _T_1017;
  assign Queue_6_io_enq_bits = io_in_0_aw_bits_user;
  assign Queue_6_io_deq_ready = _T_1015;
  assign Queue_7_clock = clock;
  assign Queue_7_reset = reset;
  assign Queue_7_io_enq_valid = _T_1021;
  assign Queue_7_io_enq_bits = io_in_0_aw_bits_user;
  assign Queue_7_io_deq_ready = _T_1019;
  assign _T_700_0 = Queue_io_enq_ready;
  assign _T_700_1 = Queue_1_io_enq_ready;
  assign _T_700_2 = Queue_2_io_enq_ready;
  assign _T_700_3 = Queue_3_io_enq_ready;
  assign _GEN_8 = 4'h1 == io_in_0_ar_bits_id ? _T_700_1 : _T_700_0;
  assign _GEN_9 = 4'h2 == io_in_0_ar_bits_id ? _T_700_2 : _GEN_8;
  assign _GEN_10 = 4'h3 == io_in_0_ar_bits_id ? _T_700_3 : _GEN_9;
  assign _GEN_11 = 4'h4 == io_in_0_ar_bits_id ? 1'h0 : _GEN_10;
  assign _GEN_12 = 4'h5 == io_in_0_ar_bits_id ? 1'h0 : _GEN_11;
  assign _GEN_13 = 4'h6 == io_in_0_ar_bits_id ? 1'h0 : _GEN_12;
  assign _GEN_14 = 4'h7 == io_in_0_ar_bits_id ? 1'h0 : _GEN_13;
  assign _GEN_15 = 4'h8 == io_in_0_ar_bits_id ? 1'h0 : _GEN_14;
  assign _GEN_16 = 4'h9 == io_in_0_ar_bits_id ? 1'h0 : _GEN_15;
  assign _GEN_17 = 4'ha == io_in_0_ar_bits_id ? 1'h0 : _GEN_16;
  assign _GEN_18 = 4'hb == io_in_0_ar_bits_id ? 1'h0 : _GEN_17;
  assign _GEN_19 = 4'hc == io_in_0_ar_bits_id ? 1'h0 : _GEN_18;
  assign _GEN_20 = 4'hd == io_in_0_ar_bits_id ? 1'h0 : _GEN_19;
  assign _GEN_21 = 4'he == io_in_0_ar_bits_id ? 1'h0 : _GEN_20;
  assign _GEN_22 = 4'hf == io_in_0_ar_bits_id ? 1'h0 : _GEN_21;
  assign _T_720 = io_out_0_ar_ready & _GEN_22;
  assign _T_721 = io_in_0_ar_valid & _GEN_22;
  assign _T_724_0 = Queue_io_deq_valid;
  assign _T_724_1 = Queue_1_io_deq_valid;
  assign _T_724_2 = Queue_2_io_deq_valid;
  assign _T_724_3 = Queue_3_io_deq_valid;
  assign _T_746_0 = Queue_io_deq_bits;
  assign _T_746_1 = Queue_1_io_deq_bits;
  assign _T_746_2 = Queue_2_io_deq_bits;
  assign _T_746_3 = Queue_3_io_deq_bits;
  assign _T_767 = io_out_0_r_valid == 1'h0;
  assign _GEN_23 = 4'h1 == io_out_0_r_bits_id ? _T_724_1 : _T_724_0;
  assign _GEN_24 = 4'h2 == io_out_0_r_bits_id ? _T_724_2 : _GEN_23;
  assign _GEN_25 = 4'h3 == io_out_0_r_bits_id ? _T_724_3 : _GEN_24;
  assign _GEN_26 = 4'h4 == io_out_0_r_bits_id ? 1'h0 : _GEN_25;
  assign _GEN_27 = 4'h5 == io_out_0_r_bits_id ? 1'h0 : _GEN_26;
  assign _GEN_28 = 4'h6 == io_out_0_r_bits_id ? 1'h0 : _GEN_27;
  assign _GEN_29 = 4'h7 == io_out_0_r_bits_id ? 1'h0 : _GEN_28;
  assign _GEN_30 = 4'h8 == io_out_0_r_bits_id ? 1'h0 : _GEN_29;
  assign _GEN_31 = 4'h9 == io_out_0_r_bits_id ? 1'h0 : _GEN_30;
  assign _GEN_32 = 4'ha == io_out_0_r_bits_id ? 1'h0 : _GEN_31;
  assign _GEN_33 = 4'hb == io_out_0_r_bits_id ? 1'h0 : _GEN_32;
  assign _GEN_34 = 4'hc == io_out_0_r_bits_id ? 1'h0 : _GEN_33;
  assign _GEN_35 = 4'hd == io_out_0_r_bits_id ? 1'h0 : _GEN_34;
  assign _GEN_36 = 4'he == io_out_0_r_bits_id ? 1'h0 : _GEN_35;
  assign _GEN_37 = 4'hf == io_out_0_r_bits_id ? 1'h0 : _GEN_36;
  assign _T_768 = _T_767 | _GEN_37;
  assign _T_769 = _T_768 | reset;
  assign _T_771 = _T_769 == 1'h0;
  assign _GEN_38 = 4'h1 == io_out_0_r_bits_id ? _T_746_1 : _T_746_0;
  assign _GEN_39 = 4'h2 == io_out_0_r_bits_id ? _T_746_2 : _GEN_38;
  assign _GEN_40 = 4'h3 == io_out_0_r_bits_id ? _T_746_3 : _GEN_39;
  assign _GEN_41 = 4'h4 == io_out_0_r_bits_id ? 12'h0 : _GEN_40;
  assign _GEN_42 = 4'h5 == io_out_0_r_bits_id ? 12'h0 : _GEN_41;
  assign _GEN_43 = 4'h6 == io_out_0_r_bits_id ? 12'h0 : _GEN_42;
  assign _GEN_44 = 4'h7 == io_out_0_r_bits_id ? 12'h0 : _GEN_43;
  assign _GEN_45 = 4'h8 == io_out_0_r_bits_id ? 12'h0 : _GEN_44;
  assign _GEN_46 = 4'h9 == io_out_0_r_bits_id ? 12'h0 : _GEN_45;
  assign _GEN_47 = 4'ha == io_out_0_r_bits_id ? 12'h0 : _GEN_46;
  assign _GEN_48 = 4'hb == io_out_0_r_bits_id ? 12'h0 : _GEN_47;
  assign _GEN_49 = 4'hc == io_out_0_r_bits_id ? 12'h0 : _GEN_48;
  assign _GEN_50 = 4'hd == io_out_0_r_bits_id ? 12'h0 : _GEN_49;
  assign _GEN_51 = 4'he == io_out_0_r_bits_id ? 12'h0 : _GEN_50;
  assign _GEN_52 = 4'hf == io_out_0_r_bits_id ? 12'h0 : _GEN_51;
  assign _T_774 = 16'h1 << io_in_0_ar_bits_id;
  assign _T_776 = _T_774[0];
  assign _T_777 = _T_774[1];
  assign _T_778 = _T_774[2];
  assign _T_779 = _T_774[3];
  assign _T_794 = 16'h1 << io_out_0_r_bits_id;
  assign _T_796 = _T_794[0];
  assign _T_797 = _T_794[1];
  assign _T_798 = _T_794[2];
  assign _T_799 = _T_794[3];
  assign _T_812 = io_out_0_r_valid & io_in_0_r_ready;
  assign _T_813 = _T_812 & _T_796;
  assign _T_814 = _T_813 & io_out_0_r_bits_last;
  assign _T_815 = io_in_0_ar_valid & io_out_0_ar_ready;
  assign _T_816 = _T_815 & _T_776;
  assign _T_818 = _T_812 & _T_797;
  assign _T_819 = _T_818 & io_out_0_r_bits_last;
  assign _T_821 = _T_815 & _T_777;
  assign _T_823 = _T_812 & _T_798;
  assign _T_824 = _T_823 & io_out_0_r_bits_last;
  assign _T_826 = _T_815 & _T_778;
  assign _T_828 = _T_812 & _T_799;
  assign _T_829 = _T_828 & io_out_0_r_bits_last;
  assign _T_831 = _T_815 & _T_779;
  assign _T_894_0 = Queue_4_io_enq_ready;
  assign _T_894_1 = Queue_5_io_enq_ready;
  assign _T_894_2 = Queue_6_io_enq_ready;
  assign _T_894_3 = Queue_7_io_enq_ready;
  assign _GEN_53 = 4'h1 == io_in_0_aw_bits_id ? _T_894_1 : _T_894_0;
  assign _GEN_54 = 4'h2 == io_in_0_aw_bits_id ? _T_894_2 : _GEN_53;
  assign _GEN_55 = 4'h3 == io_in_0_aw_bits_id ? _T_894_3 : _GEN_54;
  assign _GEN_56 = 4'h4 == io_in_0_aw_bits_id ? 1'h0 : _GEN_55;
  assign _GEN_57 = 4'h5 == io_in_0_aw_bits_id ? 1'h0 : _GEN_56;
  assign _GEN_58 = 4'h6 == io_in_0_aw_bits_id ? 1'h0 : _GEN_57;
  assign _GEN_59 = 4'h7 == io_in_0_aw_bits_id ? 1'h0 : _GEN_58;
  assign _GEN_60 = 4'h8 == io_in_0_aw_bits_id ? 1'h0 : _GEN_59;
  assign _GEN_61 = 4'h9 == io_in_0_aw_bits_id ? 1'h0 : _GEN_60;
  assign _GEN_62 = 4'ha == io_in_0_aw_bits_id ? 1'h0 : _GEN_61;
  assign _GEN_63 = 4'hb == io_in_0_aw_bits_id ? 1'h0 : _GEN_62;
  assign _GEN_64 = 4'hc == io_in_0_aw_bits_id ? 1'h0 : _GEN_63;
  assign _GEN_65 = 4'hd == io_in_0_aw_bits_id ? 1'h0 : _GEN_64;
  assign _GEN_66 = 4'he == io_in_0_aw_bits_id ? 1'h0 : _GEN_65;
  assign _GEN_67 = 4'hf == io_in_0_aw_bits_id ? 1'h0 : _GEN_66;
  assign _T_914 = io_out_0_aw_ready & _GEN_67;
  assign _T_915 = io_in_0_aw_valid & _GEN_67;
  assign _T_918_0 = Queue_4_io_deq_valid;
  assign _T_918_1 = Queue_5_io_deq_valid;
  assign _T_918_2 = Queue_6_io_deq_valid;
  assign _T_918_3 = Queue_7_io_deq_valid;
  assign _T_940_0 = Queue_4_io_deq_bits;
  assign _T_940_1 = Queue_5_io_deq_bits;
  assign _T_940_2 = Queue_6_io_deq_bits;
  assign _T_940_3 = Queue_7_io_deq_bits;
  assign _T_961 = io_out_0_b_valid == 1'h0;
  assign _GEN_68 = 4'h1 == io_out_0_b_bits_id ? _T_918_1 : _T_918_0;
  assign _GEN_69 = 4'h2 == io_out_0_b_bits_id ? _T_918_2 : _GEN_68;
  assign _GEN_70 = 4'h3 == io_out_0_b_bits_id ? _T_918_3 : _GEN_69;
  assign _GEN_71 = 4'h4 == io_out_0_b_bits_id ? 1'h0 : _GEN_70;
  assign _GEN_72 = 4'h5 == io_out_0_b_bits_id ? 1'h0 : _GEN_71;
  assign _GEN_73 = 4'h6 == io_out_0_b_bits_id ? 1'h0 : _GEN_72;
  assign _GEN_74 = 4'h7 == io_out_0_b_bits_id ? 1'h0 : _GEN_73;
  assign _GEN_75 = 4'h8 == io_out_0_b_bits_id ? 1'h0 : _GEN_74;
  assign _GEN_76 = 4'h9 == io_out_0_b_bits_id ? 1'h0 : _GEN_75;
  assign _GEN_77 = 4'ha == io_out_0_b_bits_id ? 1'h0 : _GEN_76;
  assign _GEN_78 = 4'hb == io_out_0_b_bits_id ? 1'h0 : _GEN_77;
  assign _GEN_79 = 4'hc == io_out_0_b_bits_id ? 1'h0 : _GEN_78;
  assign _GEN_80 = 4'hd == io_out_0_b_bits_id ? 1'h0 : _GEN_79;
  assign _GEN_81 = 4'he == io_out_0_b_bits_id ? 1'h0 : _GEN_80;
  assign _GEN_82 = 4'hf == io_out_0_b_bits_id ? 1'h0 : _GEN_81;
  assign _T_962 = _T_961 | _GEN_82;
  assign _T_963 = _T_962 | reset;
  assign _T_965 = _T_963 == 1'h0;
  assign _GEN_83 = 4'h1 == io_out_0_b_bits_id ? _T_940_1 : _T_940_0;
  assign _GEN_84 = 4'h2 == io_out_0_b_bits_id ? _T_940_2 : _GEN_83;
  assign _GEN_85 = 4'h3 == io_out_0_b_bits_id ? _T_940_3 : _GEN_84;
  assign _GEN_86 = 4'h4 == io_out_0_b_bits_id ? 12'h0 : _GEN_85;
  assign _GEN_87 = 4'h5 == io_out_0_b_bits_id ? 12'h0 : _GEN_86;
  assign _GEN_88 = 4'h6 == io_out_0_b_bits_id ? 12'h0 : _GEN_87;
  assign _GEN_89 = 4'h7 == io_out_0_b_bits_id ? 12'h0 : _GEN_88;
  assign _GEN_90 = 4'h8 == io_out_0_b_bits_id ? 12'h0 : _GEN_89;
  assign _GEN_91 = 4'h9 == io_out_0_b_bits_id ? 12'h0 : _GEN_90;
  assign _GEN_92 = 4'ha == io_out_0_b_bits_id ? 12'h0 : _GEN_91;
  assign _GEN_93 = 4'hb == io_out_0_b_bits_id ? 12'h0 : _GEN_92;
  assign _GEN_94 = 4'hc == io_out_0_b_bits_id ? 12'h0 : _GEN_93;
  assign _GEN_95 = 4'hd == io_out_0_b_bits_id ? 12'h0 : _GEN_94;
  assign _GEN_96 = 4'he == io_out_0_b_bits_id ? 12'h0 : _GEN_95;
  assign _GEN_97 = 4'hf == io_out_0_b_bits_id ? 12'h0 : _GEN_96;
  assign _T_968 = 16'h1 << io_in_0_aw_bits_id;
  assign _T_970 = _T_968[0];
  assign _T_971 = _T_968[1];
  assign _T_972 = _T_968[2];
  assign _T_973 = _T_968[3];
  assign _T_988 = 16'h1 << io_out_0_b_bits_id;
  assign _T_990 = _T_988[0];
  assign _T_991 = _T_988[1];
  assign _T_992 = _T_988[2];
  assign _T_993 = _T_988[3];
  assign _T_1006 = io_out_0_b_valid & io_in_0_b_ready;
  assign _T_1007 = _T_1006 & _T_990;
  assign _T_1008 = io_in_0_aw_valid & io_out_0_aw_ready;
  assign _T_1009 = _T_1008 & _T_970;
  assign _T_1011 = _T_1006 & _T_991;
  assign _T_1013 = _T_1008 & _T_971;
  assign _T_1015 = _T_1006 & _T_992;
  assign _T_1017 = _T_1008 & _T_972;
  assign _T_1019 = _T_1006 & _T_993;
  assign _T_1021 = _T_1008 & _T_973;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_771) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:60 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_771) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_965) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:81 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_965) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_25(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [30:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [30:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire  ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire  ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [30:0] ram_addr [0:1];
  reg [31:0] _RAND_1;
  wire [30:0] ram_addr__T_43_data;
  wire  ram_addr__T_43_addr;
  wire [30:0] ram_addr__T_29_data;
  wire  ram_addr__T_29_addr;
  wire  ram_addr__T_29_mask;
  wire  ram_addr__T_29_en;
  reg [7:0] ram_len [0:1];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_43_data;
  wire  ram_len__T_43_addr;
  wire [7:0] ram_len__T_29_data;
  wire  ram_len__T_29_addr;
  wire  ram_len__T_29_mask;
  wire  ram_len__T_29_en;
  reg [2:0] ram_size [0:1];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [2:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg [1:0] ram_burst [0:1];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_43_data;
  wire  ram_burst__T_43_addr;
  wire [1:0] ram_burst__T_29_data;
  wire  ram_burst__T_29_addr;
  wire  ram_burst__T_29_mask;
  wire  ram_burst__T_29_en;
  reg  value;
  reg [31:0] _RAND_5;
  reg  value_1;
  reg [31:0] _RAND_6;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_12;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_13;
  wire  _T_38;
  wire  _GEN_14;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_addr = ram_addr__T_43_data;
  assign io_deq_bits_len = ram_len__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_burst = ram_burst__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_addr__T_43_addr = value_1;
  assign ram_addr__T_43_data = ram_addr[ram_addr__T_43_addr];
  assign ram_addr__T_29_data = io_enq_bits_addr;
  assign ram_addr__T_29_addr = value;
  assign ram_addr__T_29_mask = _T_25;
  assign ram_addr__T_29_en = _T_25;
  assign ram_len__T_43_addr = value_1;
  assign ram_len__T_43_data = ram_len[ram_len__T_43_addr];
  assign ram_len__T_29_data = io_enq_bits_len;
  assign ram_len__T_29_addr = value;
  assign ram_len__T_29_mask = _T_25;
  assign ram_len__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_burst__T_43_addr = value_1;
  assign ram_burst__T_43_data = ram_burst[ram_burst__T_43_addr];
  assign ram_burst__T_29_data = io_enq_bits_burst;
  assign ram_burst__T_29_addr = value;
  assign ram_burst__T_29_mask = _T_25;
  assign ram_burst__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_12 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_13 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_14 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[30:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_addr__T_29_en & ram_addr__T_29_mask) begin
      ram_addr[ram_addr__T_29_addr] <= ram_addr__T_29_data;
    end
    if(ram_len__T_29_en & ram_len__T_29_mask) begin
      ram_len[ram_len__T_29_addr] <= ram_len__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_burst__T_29_en & ram_burst__T_29_mask) begin
      ram_burst[ram_burst__T_29_addr] <= ram_burst__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_26(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input  [7:0]  io_enq_bits_strb,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_data,
  output [7:0]  io_deq_bits_strb,
  output        io_deq_bits_last
);
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_0;
  wire [63:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [63:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] _RAND_1;
  wire [7:0] ram_strb__T_43_data;
  wire  ram_strb__T_43_addr;
  wire [7:0] ram_strb__T_29_data;
  wire  ram_strb__T_29_addr;
  wire  ram_strb__T_29_mask;
  wire  ram_strb__T_29_en;
  reg  ram_last [0:1];
  reg [31:0] _RAND_2;
  wire  ram_last__T_43_data;
  wire  ram_last__T_43_addr;
  wire  ram_last__T_29_data;
  wire  ram_last__T_29_addr;
  wire  ram_last__T_29_mask;
  wire  ram_last__T_29_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_6;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_7;
  wire  _T_38;
  wire  _GEN_8;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign io_deq_bits_strb = ram_strb__T_43_data;
  assign io_deq_bits_last = ram_last__T_43_data;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign ram_strb__T_43_addr = value_1;
  assign ram_strb__T_43_data = ram_strb[ram_strb__T_43_addr];
  assign ram_strb__T_29_data = io_enq_bits_strb;
  assign ram_strb__T_29_addr = value;
  assign ram_strb__T_29_mask = _T_25;
  assign ram_strb__T_29_en = _T_25;
  assign ram_last__T_43_addr = value_1;
  assign ram_last__T_43_data = ram_last[ram_last__T_43_addr];
  assign ram_last__T_29_data = io_enq_bits_last;
  assign ram_last__T_29_addr = value;
  assign ram_last__T_29_mask = _T_25;
  assign ram_last__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_6 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_7 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_8 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = _RAND_1[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if(ram_strb__T_29_en & ram_strb__T_29_mask) begin
      ram_strb[ram_strb__T_29_addr] <= ram_strb__T_29_data;
    end
    if(ram_last__T_29_en & ram_last__T_29_mask) begin
      ram_last[ram_last__T_29_addr] <= ram_last__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_27(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire  ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire  ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] ram_resp__T_43_data;
  wire  ram_resp__T_43_addr;
  wire [1:0] ram_resp__T_29_data;
  wire  ram_resp__T_29_addr;
  wire  ram_resp__T_29_mask;
  wire  ram_resp__T_29_en;
  reg  value;
  reg [31:0] _RAND_2;
  reg  value_1;
  reg [31:0] _RAND_3;
  reg  maybe_full;
  reg [31:0] _RAND_4;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_5;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_6;
  wire  _T_38;
  wire  _GEN_7;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_resp = ram_resp__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_resp__T_43_addr = value_1;
  assign ram_resp__T_43_data = ram_resp[ram_resp__T_43_addr];
  assign ram_resp__T_29_data = io_enq_bits_resp;
  assign ram_resp__T_29_addr = value;
  assign ram_resp__T_29_mask = _T_25;
  assign ram_resp__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_5 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_6 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_7 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  maybe_full = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_resp__T_29_en & ram_resp__T_29_mask) begin
      ram_resp[ram_resp__T_29_addr] <= ram_resp__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_29(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_last
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire  ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire  ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [63:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_43_data;
  wire  ram_resp__T_43_addr;
  wire [1:0] ram_resp__T_29_data;
  wire  ram_resp__T_29_addr;
  wire  ram_resp__T_29_mask;
  wire  ram_resp__T_29_en;
  reg  ram_last [0:1];
  reg [31:0] _RAND_3;
  wire  ram_last__T_43_data;
  wire  ram_last__T_43_addr;
  wire  ram_last__T_29_data;
  wire  ram_last__T_29_addr;
  wire  ram_last__T_29_mask;
  wire  ram_last__T_29_en;
  reg  value;
  reg [31:0] _RAND_4;
  reg  value_1;
  reg [31:0] _RAND_5;
  reg  maybe_full;
  reg [31:0] _RAND_6;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_7;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_8;
  wire  _T_38;
  wire  _GEN_9;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign io_deq_bits_resp = ram_resp__T_43_data;
  assign io_deq_bits_last = ram_last__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign ram_resp__T_43_addr = value_1;
  assign ram_resp__T_43_data = ram_resp[ram_resp__T_43_addr];
  assign ram_resp__T_29_data = io_enq_bits_resp;
  assign ram_resp__T_29_addr = value;
  assign ram_resp__T_29_mask = _T_25;
  assign ram_resp__T_29_en = _T_25;
  assign ram_last__T_43_addr = value_1;
  assign ram_last__T_43_data = ram_last[ram_last__T_43_addr];
  assign ram_last__T_29_data = io_enq_bits_last;
  assign ram_last__T_29_addr = value;
  assign ram_last__T_29_mask = _T_25;
  assign ram_last__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_7 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_8 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_9 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  maybe_full = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if(ram_resp__T_29_en & ram_resp__T_29_mask) begin
      ram_resp[ram_resp__T_29_addr] <= ram_resp__T_29_data;
    end
    if(ram_last__T_29_en & ram_last__T_29_mask) begin
      ram_last[ram_last__T_29_addr] <= ram_last__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module AXI4Buffer(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [3:0]  io_in_0_aw_bits_id,
  input  [30:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [3:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [3:0]  io_in_0_ar_bits_id,
  input  [30:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [3:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output        io_in_0_r_bits_last,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [3:0]  io_out_0_aw_bits_id,
  output [30:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [1:0]  io_out_0_aw_bits_burst,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [3:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [3:0]  io_out_0_ar_bits_id,
  output [30:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [1:0]  io_out_0_ar_bits_burst,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [3:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input         io_out_0_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [30:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [30:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire  _T_95_valid;
  wire [3:0] _T_95_bits_id;
  wire [30:0] _T_95_bits_addr;
  wire [7:0] _T_95_bits_len;
  wire [2:0] _T_95_bits_size;
  wire [1:0] _T_95_bits_burst;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [7:0] Queue_1_io_enq_bits_strb;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [7:0] Queue_1_io_deq_bits_strb;
  wire  Queue_1_io_deq_bits_last;
  wire  _T_104_valid;
  wire [63:0] _T_104_bits_data;
  wire [7:0] _T_104_bits_strb;
  wire  _T_104_bits_last;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire  _T_113_valid;
  wire [3:0] _T_113_bits_id;
  wire [1:0] _T_113_bits_resp;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [30:0] Queue_3_io_enq_bits_addr;
  wire [7:0] Queue_3_io_enq_bits_len;
  wire [2:0] Queue_3_io_enq_bits_size;
  wire [1:0] Queue_3_io_enq_bits_burst;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [30:0] Queue_3_io_deq_bits_addr;
  wire [7:0] Queue_3_io_deq_bits_len;
  wire [2:0] Queue_3_io_deq_bits_size;
  wire [1:0] Queue_3_io_deq_bits_burst;
  wire  _T_122_valid;
  wire [3:0] _T_122_bits_id;
  wire [30:0] _T_122_bits_addr;
  wire [7:0] _T_122_bits_len;
  wire [2:0] _T_122_bits_size;
  wire [1:0] _T_122_bits_burst;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire  Queue_4_io_enq_bits_last;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire  Queue_4_io_deq_bits_last;
  wire  _T_131_valid;
  wire [3:0] _T_131_bits_id;
  wire [63:0] _T_131_bits_data;
  wire [1:0] _T_131_bits_resp;
  wire  _T_131_bits_last;
  Queue_25 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst)
  );
  Queue_26 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_27 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp)
  );
  Queue_25 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_len(Queue_3_io_enq_bits_len),
    .io_enq_bits_size(Queue_3_io_enq_bits_size),
    .io_enq_bits_burst(Queue_3_io_enq_bits_burst),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_len(Queue_3_io_deq_bits_len),
    .io_deq_bits_size(Queue_3_io_deq_bits_size),
    .io_deq_bits_burst(Queue_3_io_deq_bits_burst)
  );
  Queue_29 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign io_in_0_aw_ready = Queue_io_enq_ready;
  assign io_in_0_w_ready = Queue_1_io_enq_ready;
  assign io_in_0_b_valid = _T_113_valid;
  assign io_in_0_b_bits_id = _T_113_bits_id;
  assign io_in_0_b_bits_resp = _T_113_bits_resp;
  assign io_in_0_ar_ready = Queue_3_io_enq_ready;
  assign io_in_0_r_valid = _T_131_valid;
  assign io_in_0_r_bits_id = _T_131_bits_id;
  assign io_in_0_r_bits_data = _T_131_bits_data;
  assign io_in_0_r_bits_resp = _T_131_bits_resp;
  assign io_in_0_r_bits_last = _T_131_bits_last;
  assign io_out_0_aw_valid = _T_95_valid;
  assign io_out_0_aw_bits_id = _T_95_bits_id;
  assign io_out_0_aw_bits_addr = _T_95_bits_addr;
  assign io_out_0_aw_bits_len = _T_95_bits_len;
  assign io_out_0_aw_bits_size = _T_95_bits_size;
  assign io_out_0_aw_bits_burst = _T_95_bits_burst;
  assign io_out_0_w_valid = _T_104_valid;
  assign io_out_0_w_bits_data = _T_104_bits_data;
  assign io_out_0_w_bits_strb = _T_104_bits_strb;
  assign io_out_0_w_bits_last = _T_104_bits_last;
  assign io_out_0_b_ready = Queue_2_io_enq_ready;
  assign io_out_0_ar_valid = _T_122_valid;
  assign io_out_0_ar_bits_id = _T_122_bits_id;
  assign io_out_0_ar_bits_addr = _T_122_bits_addr;
  assign io_out_0_ar_bits_len = _T_122_bits_len;
  assign io_out_0_ar_bits_size = _T_122_bits_size;
  assign io_out_0_ar_bits_burst = _T_122_bits_burst;
  assign io_out_0_r_ready = Queue_4_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_aw_valid;
  assign Queue_io_enq_bits_id = io_in_0_aw_bits_id;
  assign Queue_io_enq_bits_addr = io_in_0_aw_bits_addr;
  assign Queue_io_enq_bits_len = io_in_0_aw_bits_len;
  assign Queue_io_enq_bits_size = io_in_0_aw_bits_size;
  assign Queue_io_enq_bits_burst = io_in_0_aw_bits_burst;
  assign Queue_io_deq_ready = io_out_0_aw_ready;
  assign _T_95_valid = Queue_io_deq_valid;
  assign _T_95_bits_id = Queue_io_deq_bits_id;
  assign _T_95_bits_addr = Queue_io_deq_bits_addr;
  assign _T_95_bits_len = Queue_io_deq_bits_len;
  assign _T_95_bits_size = Queue_io_deq_bits_size;
  assign _T_95_bits_burst = Queue_io_deq_bits_burst;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_in_0_w_valid;
  assign Queue_1_io_enq_bits_data = io_in_0_w_bits_data;
  assign Queue_1_io_enq_bits_strb = io_in_0_w_bits_strb;
  assign Queue_1_io_enq_bits_last = io_in_0_w_bits_last;
  assign Queue_1_io_deq_ready = io_out_0_w_ready;
  assign _T_104_valid = Queue_1_io_deq_valid;
  assign _T_104_bits_data = Queue_1_io_deq_bits_data;
  assign _T_104_bits_strb = Queue_1_io_deq_bits_strb;
  assign _T_104_bits_last = Queue_1_io_deq_bits_last;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = io_out_0_b_valid;
  assign Queue_2_io_enq_bits_id = io_out_0_b_bits_id;
  assign Queue_2_io_enq_bits_resp = io_out_0_b_bits_resp;
  assign Queue_2_io_deq_ready = io_in_0_b_ready;
  assign _T_113_valid = Queue_2_io_deq_valid;
  assign _T_113_bits_id = Queue_2_io_deq_bits_id;
  assign _T_113_bits_resp = Queue_2_io_deq_bits_resp;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = io_in_0_ar_valid;
  assign Queue_3_io_enq_bits_id = io_in_0_ar_bits_id;
  assign Queue_3_io_enq_bits_addr = io_in_0_ar_bits_addr;
  assign Queue_3_io_enq_bits_len = io_in_0_ar_bits_len;
  assign Queue_3_io_enq_bits_size = io_in_0_ar_bits_size;
  assign Queue_3_io_enq_bits_burst = io_in_0_ar_bits_burst;
  assign Queue_3_io_deq_ready = io_out_0_ar_ready;
  assign _T_122_valid = Queue_3_io_deq_valid;
  assign _T_122_bits_id = Queue_3_io_deq_bits_id;
  assign _T_122_bits_addr = Queue_3_io_deq_bits_addr;
  assign _T_122_bits_len = Queue_3_io_deq_bits_len;
  assign _T_122_bits_size = Queue_3_io_deq_bits_size;
  assign _T_122_bits_burst = Queue_3_io_deq_bits_burst;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = io_out_0_r_valid;
  assign Queue_4_io_enq_bits_id = io_out_0_r_bits_id;
  assign Queue_4_io_enq_bits_data = io_out_0_r_bits_data;
  assign Queue_4_io_enq_bits_resp = io_out_0_r_bits_resp;
  assign Queue_4_io_enq_bits_last = io_out_0_r_bits_last;
  assign Queue_4_io_deq_ready = io_in_0_r_ready;
  assign _T_131_valid = Queue_4_io_deq_valid;
  assign _T_131_bits_id = Queue_4_io_deq_bits_id;
  assign _T_131_bits_data = Queue_4_io_deq_bits_data;
  assign _T_131_bits_resp = Queue_4_io_deq_bits_resp;
  assign _T_131_bits_last = Queue_4_io_deq_bits_last;
endmodule
module Queue_30(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [3:0]  io_enq_bits_mask,
  input  [31:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [3:0]  io_deq_bits_mask,
  output [31:0] io_deq_bits_data
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_43_data;
  wire  ram_opcode__T_43_addr;
  wire [2:0] ram_opcode__T_29_data;
  wire  ram_opcode__T_29_addr;
  wire  ram_opcode__T_29_mask;
  wire  ram_opcode__T_29_en;
  reg [2:0] ram_param [0:1];
  reg [31:0] _RAND_1;
  wire [2:0] ram_param__T_43_data;
  wire  ram_param__T_43_addr;
  wire [2:0] ram_param__T_29_data;
  wire  ram_param__T_29_addr;
  wire  ram_param__T_29_mask;
  wire  ram_param__T_29_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [3:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg [3:0] ram_source [0:1];
  reg [31:0] _RAND_3;
  wire [3:0] ram_source__T_43_data;
  wire  ram_source__T_43_addr;
  wire [3:0] ram_source__T_29_data;
  wire  ram_source__T_29_addr;
  wire  ram_source__T_29_mask;
  wire  ram_source__T_29_en;
  reg [31:0] ram_address [0:1];
  reg [31:0] _RAND_4;
  wire [31:0] ram_address__T_43_data;
  wire  ram_address__T_43_addr;
  wire [31:0] ram_address__T_29_data;
  wire  ram_address__T_29_addr;
  wire  ram_address__T_29_mask;
  wire  ram_address__T_29_en;
  reg [3:0] ram_mask [0:1];
  reg [31:0] _RAND_5;
  wire [3:0] ram_mask__T_43_data;
  wire  ram_mask__T_43_addr;
  wire [3:0] ram_mask__T_29_data;
  wire  ram_mask__T_29_addr;
  wire  ram_mask__T_29_mask;
  wire  ram_mask__T_29_en;
  reg [31:0] ram_data [0:1];
  reg [31:0] _RAND_6;
  wire [31:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [31:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg  value;
  reg [31:0] _RAND_7;
  reg  value_1;
  reg [31:0] _RAND_8;
  reg  maybe_full;
  reg [31:0] _RAND_9;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_10;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_11;
  wire  _T_38;
  wire  _GEN_12;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_opcode = ram_opcode__T_43_data;
  assign io_deq_bits_param = ram_param__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_source = ram_source__T_43_data;
  assign io_deq_bits_address = ram_address__T_43_data;
  assign io_deq_bits_mask = ram_mask__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign ram_opcode__T_43_addr = value_1;
  assign ram_opcode__T_43_data = ram_opcode[ram_opcode__T_43_addr];
  assign ram_opcode__T_29_data = io_enq_bits_opcode;
  assign ram_opcode__T_29_addr = value;
  assign ram_opcode__T_29_mask = _T_25;
  assign ram_opcode__T_29_en = _T_25;
  assign ram_param__T_43_addr = value_1;
  assign ram_param__T_43_data = ram_param[ram_param__T_43_addr];
  assign ram_param__T_29_data = io_enq_bits_param;
  assign ram_param__T_29_addr = value;
  assign ram_param__T_29_mask = _T_25;
  assign ram_param__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_source__T_43_addr = value_1;
  assign ram_source__T_43_data = ram_source[ram_source__T_43_addr];
  assign ram_source__T_29_data = io_enq_bits_source;
  assign ram_source__T_29_addr = value;
  assign ram_source__T_29_mask = _T_25;
  assign ram_source__T_29_en = _T_25;
  assign ram_address__T_43_addr = value_1;
  assign ram_address__T_43_data = ram_address[ram_address__T_43_addr];
  assign ram_address__T_29_data = io_enq_bits_address;
  assign ram_address__T_29_addr = value;
  assign ram_address__T_29_mask = _T_25;
  assign ram_address__T_29_en = _T_25;
  assign ram_mask__T_43_addr = value_1;
  assign ram_mask__T_43_data = ram_mask[ram_mask__T_43_addr];
  assign ram_mask__T_29_data = io_enq_bits_mask;
  assign ram_mask__T_29_addr = value;
  assign ram_mask__T_29_mask = _T_25;
  assign ram_mask__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_10 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_11 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_12 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_address[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_mask[initvar] = _RAND_5[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  value = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  value_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  maybe_full = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_29_en & ram_opcode__T_29_mask) begin
      ram_opcode[ram_opcode__T_29_addr] <= ram_opcode__T_29_data;
    end
    if(ram_param__T_29_en & ram_param__T_29_mask) begin
      ram_param[ram_param__T_29_addr] <= ram_param__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_source__T_29_en & ram_source__T_29_mask) begin
      ram_source[ram_source__T_29_addr] <= ram_source__T_29_data;
    end
    if(ram_address__T_29_en & ram_address__T_29_mask) begin
      ram_address[ram_address__T_29_addr] <= ram_address__T_29_data;
    end
    if(ram_mask__T_29_en & ram_mask__T_29_mask) begin
      ram_mask[ram_mask__T_29_addr] <= ram_mask__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_31(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [3:0] io_enq_bits_size,
  input  [3:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [3:0] io_deq_bits_size,
  output [3:0] io_deq_bits_source
);
  reg [2:0] ram_opcode [0:1];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_43_data;
  wire  ram_opcode__T_43_addr;
  wire [2:0] ram_opcode__T_29_data;
  wire  ram_opcode__T_29_addr;
  wire  ram_opcode__T_29_mask;
  wire  ram_opcode__T_29_en;
  reg [3:0] ram_size [0:1];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_43_data;
  wire  ram_size__T_43_addr;
  wire [3:0] ram_size__T_29_data;
  wire  ram_size__T_29_addr;
  wire  ram_size__T_29_mask;
  wire  ram_size__T_29_en;
  reg [3:0] ram_source [0:1];
  reg [31:0] _RAND_2;
  wire [3:0] ram_source__T_43_data;
  wire  ram_source__T_43_addr;
  wire [3:0] ram_source__T_29_data;
  wire  ram_source__T_29_addr;
  wire  ram_source__T_29_mask;
  wire  ram_source__T_29_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_10;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_11;
  wire  _T_38;
  wire  _GEN_12;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_opcode = ram_opcode__T_43_data;
  assign io_deq_bits_size = ram_size__T_43_data;
  assign io_deq_bits_source = ram_source__T_43_data;
  assign ram_opcode__T_43_addr = value_1;
  assign ram_opcode__T_43_data = ram_opcode[ram_opcode__T_43_addr];
  assign ram_opcode__T_29_data = io_enq_bits_opcode;
  assign ram_opcode__T_29_addr = value;
  assign ram_opcode__T_29_mask = _T_25;
  assign ram_opcode__T_29_en = _T_25;
  assign ram_size__T_43_addr = value_1;
  assign ram_size__T_43_data = ram_size[ram_size__T_43_addr];
  assign ram_size__T_29_data = io_enq_bits_size;
  assign ram_size__T_29_addr = value;
  assign ram_size__T_29_mask = _T_25;
  assign ram_size__T_29_en = _T_25;
  assign ram_source__T_43_addr = value_1;
  assign ram_source__T_43_data = ram_source[ram_source__T_43_addr];
  assign ram_source__T_29_data = io_enq_bits_source;
  assign ram_source__T_29_addr = value;
  assign ram_source__T_29_mask = _T_25;
  assign ram_source__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_10 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_11 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_12 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_29_en & ram_opcode__T_29_mask) begin
      ram_opcode[ram_opcode__T_29_addr] <= ram_opcode__T_29_data;
    end
    if(ram_size__T_29_en & ram_size__T_29_mask) begin
      ram_size[ram_size__T_29_addr] <= ram_size__T_29_data;
    end
    if(ram_source__T_29_en & ram_source__T_29_mask) begin
      ram_source[ram_source__T_29_addr] <= ram_source__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module TLBuffer_5(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input  [3:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [3:0]  io_in_0_a_bits_mask,
  input  [31:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output [3:0]  io_in_0_d_bits_source,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output [3:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input  [3:0]  io_out_0_d_bits_source
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [2:0] Queue_io_enq_bits_param;
  wire [3:0] Queue_io_enq_bits_size;
  wire [3:0] Queue_io_enq_bits_source;
  wire [31:0] Queue_io_enq_bits_address;
  wire [3:0] Queue_io_enq_bits_mask;
  wire [31:0] Queue_io_enq_bits_data;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [2:0] Queue_io_deq_bits_param;
  wire [3:0] Queue_io_deq_bits_size;
  wire [3:0] Queue_io_deq_bits_source;
  wire [31:0] Queue_io_deq_bits_address;
  wire [3:0] Queue_io_deq_bits_mask;
  wire [31:0] Queue_io_deq_bits_data;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [3:0] Queue_1_io_enq_bits_size;
  wire [3:0] Queue_1_io_enq_bits_source;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [3:0] Queue_1_io_deq_bits_size;
  wire [3:0] Queue_1_io_deq_bits_source;
  Queue_30 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_io_enq_bits_param),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_enq_bits_address(Queue_io_enq_bits_address),
    .io_enq_bits_mask(Queue_io_enq_bits_mask),
    .io_enq_bits_data(Queue_io_enq_bits_data),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_io_deq_bits_param),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source),
    .io_deq_bits_address(Queue_io_deq_bits_address),
    .io_deq_bits_mask(Queue_io_deq_bits_mask),
    .io_deq_bits_data(Queue_io_deq_bits_data)
  );
  Queue_31 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source)
  );
  assign io_in_0_a_ready = Queue_io_enq_ready;
  assign io_in_0_d_valid = Queue_1_io_deq_valid;
  assign io_in_0_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign io_in_0_d_bits_size = Queue_1_io_deq_bits_size;
  assign io_in_0_d_bits_source = Queue_1_io_deq_bits_source;
  assign io_out_0_a_valid = Queue_io_deq_valid;
  assign io_out_0_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign io_out_0_a_bits_param = Queue_io_deq_bits_param;
  assign io_out_0_a_bits_size = Queue_io_deq_bits_size;
  assign io_out_0_a_bits_source = Queue_io_deq_bits_source;
  assign io_out_0_a_bits_address = Queue_io_deq_bits_address;
  assign io_out_0_a_bits_mask = Queue_io_deq_bits_mask;
  assign io_out_0_a_bits_data = Queue_io_deq_bits_data;
  assign io_out_0_d_ready = Queue_1_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_a_valid;
  assign Queue_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Queue_io_enq_bits_param = io_in_0_a_bits_param;
  assign Queue_io_enq_bits_size = io_in_0_a_bits_size;
  assign Queue_io_enq_bits_source = io_in_0_a_bits_source;
  assign Queue_io_enq_bits_address = io_in_0_a_bits_address;
  assign Queue_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Queue_io_enq_bits_data = io_in_0_a_bits_data;
  assign Queue_io_deq_ready = io_out_0_a_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_out_0_d_valid;
  assign Queue_1_io_enq_bits_opcode = io_out_0_d_bits_opcode;
  assign Queue_1_io_enq_bits_size = io_out_0_d_bits_size;
  assign Queue_1_io_enq_bits_source = io_out_0_d_bits_source;
  assign Queue_1_io_deq_ready = io_in_0_d_ready;
endmodule
module AXI4IdIndexer_1(
  input         io_in_0_aw_valid,
  input  [7:0]  io_in_0_aw_bits_id,
  input  [31:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  input         io_in_0_ar_valid,
  input  [7:0]  io_in_0_ar_bits_id,
  input  [31:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input         io_in_0_r_ready,
  output        io_out_0_aw_valid,
  output        io_out_0_aw_bits_id,
  output [31:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [1:0]  io_out_0_aw_bits_burst,
  output [6:0]  io_out_0_aw_bits_user,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  output        io_out_0_ar_valid,
  output        io_out_0_ar_bits_id,
  output [31:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [1:0]  io_out_0_ar_bits_burst,
  output [6:0]  io_out_0_ar_bits_user,
  output        io_out_0_r_ready
);
  wire [6:0] _T_90;
  wire [6:0] _T_91;
  assign io_out_0_aw_valid = io_in_0_aw_valid;
  assign io_out_0_aw_bits_id = io_in_0_aw_bits_id[0];
  assign io_out_0_aw_bits_addr = io_in_0_aw_bits_addr;
  assign io_out_0_aw_bits_len = io_in_0_aw_bits_len;
  assign io_out_0_aw_bits_size = io_in_0_aw_bits_size;
  assign io_out_0_aw_bits_burst = io_in_0_aw_bits_burst;
  assign io_out_0_aw_bits_user = _T_91;
  assign io_out_0_w_valid = io_in_0_w_valid;
  assign io_out_0_w_bits_data = io_in_0_w_bits_data;
  assign io_out_0_w_bits_strb = io_in_0_w_bits_strb;
  assign io_out_0_w_bits_last = io_in_0_w_bits_last;
  assign io_out_0_b_ready = io_in_0_b_ready;
  assign io_out_0_ar_valid = io_in_0_ar_valid;
  assign io_out_0_ar_bits_id = io_in_0_ar_bits_id[0];
  assign io_out_0_ar_bits_addr = io_in_0_ar_bits_addr;
  assign io_out_0_ar_bits_len = io_in_0_ar_bits_len;
  assign io_out_0_ar_bits_size = io_in_0_ar_bits_size;
  assign io_out_0_ar_bits_burst = io_in_0_ar_bits_burst;
  assign io_out_0_ar_bits_user = _T_90;
  assign io_out_0_r_ready = io_in_0_r_ready;
  assign _T_90 = io_in_0_ar_bits_id[7:1];
  assign _T_91 = io_in_0_aw_bits_id[7:1];
endmodule
module Queue_32(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits_id,
  input  [31:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input  [6:0]  io_enq_bits_user,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_id,
  output [31:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst,
  output [6:0]  io_deq_bits_user
);
  reg  ram_id [0:0];
  reg [31:0] _RAND_0;
  wire  ram_id__T_35_data;
  wire  ram_id__T_35_addr;
  wire  ram_id__T_26_data;
  wire  ram_id__T_26_addr;
  wire  ram_id__T_26_mask;
  wire  ram_id__T_26_en;
  reg [31:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [31:0] ram_addr__T_35_data;
  wire  ram_addr__T_35_addr;
  wire [31:0] ram_addr__T_26_data;
  wire  ram_addr__T_26_addr;
  wire  ram_addr__T_26_mask;
  wire  ram_addr__T_26_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_35_data;
  wire  ram_len__T_35_addr;
  wire [7:0] ram_len__T_26_data;
  wire  ram_len__T_26_addr;
  wire  ram_len__T_26_mask;
  wire  ram_len__T_26_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [2:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_35_data;
  wire  ram_burst__T_35_addr;
  wire [1:0] ram_burst__T_26_data;
  wire  ram_burst__T_26_addr;
  wire  ram_burst__T_26_mask;
  wire  ram_burst__T_26_en;
  reg [6:0] ram_user [0:0];
  reg [31:0] _RAND_5;
  wire [6:0] ram_user__T_35_data;
  wire  ram_user__T_35_addr;
  wire [6:0] ram_user__T_26_data;
  wire  ram_user__T_26_addr;
  wire  ram_user__T_26_mask;
  wire  ram_user__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_6;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_13;
  wire  _T_31;
  wire  _GEN_14;
  wire  _GEN_15;
  wire  _GEN_16;
  wire [31:0] _GEN_17;
  wire [7:0] _GEN_18;
  wire [2:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [6:0] _GEN_25;
  wire  _GEN_26;
  wire  _GEN_27;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_14;
  assign io_deq_bits_id = _GEN_16;
  assign io_deq_bits_addr = _GEN_17;
  assign io_deq_bits_len = _GEN_18;
  assign io_deq_bits_size = _GEN_19;
  assign io_deq_bits_burst = _GEN_20;
  assign io_deq_bits_user = _GEN_25;
  assign ram_id__T_35_addr = 1'h0;
  assign ram_id__T_35_data = ram_id[ram_id__T_35_addr];
  assign ram_id__T_26_data = io_enq_bits_id;
  assign ram_id__T_26_addr = 1'h0;
  assign ram_id__T_26_mask = _GEN_27;
  assign ram_id__T_26_en = _GEN_27;
  assign ram_addr__T_35_addr = 1'h0;
  assign ram_addr__T_35_data = ram_addr[ram_addr__T_35_addr];
  assign ram_addr__T_26_data = io_enq_bits_addr;
  assign ram_addr__T_26_addr = 1'h0;
  assign ram_addr__T_26_mask = _GEN_27;
  assign ram_addr__T_26_en = _GEN_27;
  assign ram_len__T_35_addr = 1'h0;
  assign ram_len__T_35_data = ram_len[ram_len__T_35_addr];
  assign ram_len__T_26_data = io_enq_bits_len;
  assign ram_len__T_26_addr = 1'h0;
  assign ram_len__T_26_mask = _GEN_27;
  assign ram_len__T_26_en = _GEN_27;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_27;
  assign ram_size__T_26_en = _GEN_27;
  assign ram_burst__T_35_addr = 1'h0;
  assign ram_burst__T_35_data = ram_burst[ram_burst__T_35_addr];
  assign ram_burst__T_26_data = io_enq_bits_burst;
  assign ram_burst__T_26_addr = 1'h0;
  assign ram_burst__T_26_mask = _GEN_27;
  assign ram_burst__T_26_en = _GEN_27;
  assign ram_user__T_35_addr = 1'h0;
  assign ram_user__T_35_data = ram_user[ram_user__T_35_addr];
  assign ram_user__T_26_data = io_enq_bits_user;
  assign ram_user__T_26_addr = 1'h0;
  assign ram_user__T_26_mask = _GEN_27;
  assign ram_user__T_26_en = _GEN_27;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_27 != _GEN_26;
  assign _GEN_13 = _T_29 ? _GEN_27 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_14 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_15 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_16 = _T_18 ? io_enq_bits_id : ram_id__T_35_data;
  assign _GEN_17 = _T_18 ? io_enq_bits_addr : ram_addr__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_len : ram_len__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_20 = _T_18 ? io_enq_bits_burst : ram_burst__T_35_data;
  assign _GEN_25 = _T_18 ? io_enq_bits_user : ram_user__T_35_data;
  assign _GEN_26 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_27 = _T_18 ? _GEN_15 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = _RAND_5[6:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  maybe_full = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_26_en & ram_id__T_26_mask) begin
      ram_id[ram_id__T_26_addr] <= ram_id__T_26_data;
    end
    if(ram_addr__T_26_en & ram_addr__T_26_mask) begin
      ram_addr[ram_addr__T_26_addr] <= ram_addr__T_26_data;
    end
    if(ram_len__T_26_en & ram_len__T_26_mask) begin
      ram_len[ram_len__T_26_addr] <= ram_len__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_burst__T_26_en & ram_burst__T_26_mask) begin
      ram_burst[ram_burst__T_26_addr] <= ram_burst__T_26_data;
    end
    if(ram_user__T_26_en & ram_user__T_26_mask) begin
      ram_user[ram_user__T_26_addr] <= ram_user__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module AXI4Fragmenter(
  input         clock,
  input         reset,
  input         io_in_0_aw_valid,
  input         io_in_0_aw_bits_id,
  input  [31:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  input  [6:0]  io_in_0_aw_bits_user,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  input         io_in_0_ar_valid,
  input         io_in_0_ar_bits_id,
  input  [31:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input  [6:0]  io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output        io_out_0_aw_bits_id,
  output [31:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  output [7:0]  io_out_0_aw_bits_user,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input  [7:0]  io_out_0_b_bits_user,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output        io_out_0_ar_bits_id,
  output [31:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output [7:0]  io_out_0_ar_bits_user,
  output        io_out_0_r_ready
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire  Queue_io_enq_bits_id;
  wire [31:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire [6:0] Queue_io_enq_bits_user;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire  Queue_io_deq_bits_id;
  wire [31:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire [6:0] Queue_io_deq_bits_user;
  wire  _T_95_valid;
  wire  _T_95_bits_id;
  wire [31:0] _T_95_bits_addr;
  wire [7:0] _T_95_bits_len;
  wire [2:0] _T_95_bits_size;
  wire [1:0] _T_95_bits_burst;
  wire [6:0] _T_95_bits_user;
  reg  _T_105;
  reg [31:0] _RAND_0;
  reg [31:0] _T_107;
  reg [31:0] _RAND_1;
  reg [7:0] _T_109;
  reg [31:0] _RAND_2;
  wire [7:0] _T_110;
  wire [31:0] _T_111;
  wire [28:0] _T_113;
  wire [7:0] _T_114;
  wire [31:0] _T_116;
  wire [32:0] _T_117;
  wire [32:0] _T_119;
  wire [32:0] _T_120;
  wire  _T_122;
  wire [31:0] _T_124;
  wire [32:0] _T_125;
  wire [32:0] _T_127;
  wire [32:0] _T_128;
  wire  _T_130;
  wire [32:0] _T_133;
  wire [32:0] _T_135;
  wire [32:0] _T_136;
  wire  _T_138;
  wire [31:0] _T_140;
  wire [32:0] _T_141;
  wire [32:0] _T_143;
  wire [32:0] _T_144;
  wire  _T_146;
  wire [31:0] _T_148;
  wire [32:0] _T_149;
  wire [32:0] _T_151;
  wire [32:0] _T_152;
  wire  _T_154;
  wire [31:0] _T_156;
  wire [32:0] _T_157;
  wire [32:0] _T_159;
  wire [32:0] _T_160;
  wire  _T_162;
  wire  _T_163;
  wire  _T_164;
  wire  _T_165;
  wire  _T_166;
  wire  _T_167;
  wire [31:0] _T_170;
  wire [32:0] _T_171;
  wire [32:0] _T_173;
  wire [32:0] _T_174;
  wire  _T_176;
  wire [2:0] _T_180;
  wire [7:0] _T_182;
  wire [7:0] _GEN_16;
  wire [7:0] _T_183;
  wire [6:0] _T_186;
  wire [7:0] _GEN_17;
  wire [7:0] _T_187;
  wire [5:0] _T_188;
  wire [7:0] _GEN_18;
  wire [7:0] _T_189;
  wire [3:0] _T_190;
  wire [7:0] _GEN_19;
  wire [7:0] _T_191;
  wire [6:0] _T_193;
  wire [7:0] _T_194;
  wire [8:0] _GEN_20;
  wire [8:0] _T_195;
  wire [7:0] _T_196;
  wire [7:0] _T_197;
  wire [9:0] _GEN_21;
  wire [9:0] _T_198;
  wire [7:0] _T_199;
  wire [7:0] _T_200;
  wire [11:0] _GEN_22;
  wire [11:0] _T_201;
  wire [7:0] _T_202;
  wire [7:0] _T_203;
  wire [7:0] _T_205;
  wire [7:0] _GEN_23;
  wire [7:0] _T_206;
  wire [8:0] _GEN_24;
  wire [8:0] _T_207;
  wire [7:0] _T_208;
  wire [7:0] _T_209;
  wire [9:0] _GEN_25;
  wire [9:0] _T_210;
  wire [7:0] _T_211;
  wire [7:0] _T_212;
  wire [11:0] _GEN_26;
  wire [11:0] _T_213;
  wire [7:0] _T_214;
  wire [7:0] _T_215;
  wire [7:0] _T_217;
  wire [7:0] _T_218;
  wire [7:0] _T_219;
  wire  _T_221;
  wire  _T_223;
  wire  _T_224;
  wire [7:0] _T_226;
  wire [8:0] _GEN_27;
  wire [8:0] _T_227;
  wire [8:0] _T_229;
  wire [8:0] _T_231;
  wire [8:0] _T_232;
  wire [8:0] _T_233;
  wire [15:0] _GEN_28;
  wire [15:0] _T_234;
  wire [31:0] _GEN_29;
  wire [32:0] _T_235;
  wire [31:0] _T_236;
  wire [15:0] _T_238;
  wire [22:0] _GEN_30;
  wire [22:0] _T_239;
  wire [14:0] _T_240;
  wire  _T_244;
  wire [31:0] _GEN_31;
  wire [31:0] _T_245;
  wire [31:0] _T_246;
  wire [31:0] _T_247;
  wire [31:0] _T_248;
  wire [31:0] _T_249;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire  _T_252;
  wire  _T_253;
  wire [31:0] _T_254;
  wire [9:0] _T_257;
  wire [2:0] _T_258;
  wire [2:0] _T_259;
  wire [31:0] _GEN_33;
  wire [31:0] _T_260;
  wire [31:0] _T_261;
  wire  _T_262;
  wire  _T_264;
  wire [8:0] _GEN_34;
  wire [9:0] _T_265;
  wire [9:0] _T_266;
  wire [8:0] _T_267;
  wire  _GEN_3;
  wire [31:0] _GEN_4;
  wire [8:0] _GEN_5;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire  Queue_1_io_enq_bits_id;
  wire [31:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [1:0] Queue_1_io_enq_bits_burst;
  wire [6:0] Queue_1_io_enq_bits_user;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire  Queue_1_io_deq_bits_id;
  wire [31:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire [6:0] Queue_1_io_deq_bits_user;
  wire  _T_273_valid;
  wire  _T_273_bits_id;
  wire [31:0] _T_273_bits_addr;
  wire [7:0] _T_273_bits_len;
  wire [2:0] _T_273_bits_size;
  wire [1:0] _T_273_bits_burst;
  wire [6:0] _T_273_bits_user;
  reg  _T_283;
  reg [31:0] _RAND_3;
  reg [31:0] _T_285;
  reg [31:0] _RAND_4;
  reg [7:0] _T_287;
  reg [31:0] _RAND_5;
  wire [7:0] _T_288;
  wire [31:0] _T_289;
  wire [28:0] _T_291;
  wire [7:0] _T_292;
  wire [31:0] _T_294;
  wire [32:0] _T_295;
  wire [32:0] _T_297;
  wire [32:0] _T_298;
  wire  _T_300;
  wire [31:0] _T_303;
  wire [32:0] _T_304;
  wire [32:0] _T_306;
  wire [32:0] _T_307;
  wire  _T_309;
  wire [31:0] _T_311;
  wire [32:0] _T_312;
  wire [32:0] _T_314;
  wire [32:0] _T_315;
  wire  _T_317;
  wire [32:0] _T_320;
  wire [32:0] _T_322;
  wire [32:0] _T_323;
  wire  _T_325;
  wire [31:0] _T_327;
  wire [32:0] _T_328;
  wire [32:0] _T_330;
  wire [32:0] _T_331;
  wire  _T_333;
  wire  _T_334;
  wire  _T_335;
  wire  _T_336;
  wire [31:0] _T_339;
  wire [32:0] _T_340;
  wire [32:0] _T_342;
  wire [32:0] _T_343;
  wire  _T_345;
  wire [4:0] _T_349;
  wire [2:0] _T_351;
  wire [7:0] _T_353;
  wire [4:0] _GEN_35;
  wire [4:0] _T_354;
  wire [7:0] _GEN_36;
  wire [7:0] _T_355;
  wire [6:0] _T_358;
  wire [7:0] _GEN_37;
  wire [7:0] _T_359;
  wire [5:0] _T_360;
  wire [7:0] _GEN_38;
  wire [7:0] _T_361;
  wire [3:0] _T_362;
  wire [7:0] _GEN_39;
  wire [7:0] _T_363;
  wire [6:0] _T_365;
  wire [7:0] _T_366;
  wire [8:0] _GEN_40;
  wire [8:0] _T_367;
  wire [7:0] _T_368;
  wire [7:0] _T_369;
  wire [9:0] _GEN_41;
  wire [9:0] _T_370;
  wire [7:0] _T_371;
  wire [7:0] _T_372;
  wire [11:0] _GEN_42;
  wire [11:0] _T_373;
  wire [7:0] _T_374;
  wire [7:0] _T_375;
  wire [7:0] _T_377;
  wire [7:0] _GEN_43;
  wire [7:0] _T_378;
  wire [8:0] _GEN_44;
  wire [8:0] _T_379;
  wire [7:0] _T_380;
  wire [7:0] _T_381;
  wire [9:0] _GEN_45;
  wire [9:0] _T_382;
  wire [7:0] _T_383;
  wire [7:0] _T_384;
  wire [11:0] _GEN_46;
  wire [11:0] _T_385;
  wire [7:0] _T_386;
  wire [7:0] _T_387;
  wire [7:0] _T_389;
  wire [7:0] _T_390;
  wire [7:0] _T_391;
  wire  _T_393;
  wire  _T_395;
  wire  _T_396;
  wire [7:0] _T_398;
  wire [8:0] _GEN_47;
  wire [8:0] _T_399;
  wire [8:0] _T_401;
  wire [8:0] _T_403;
  wire [8:0] _T_404;
  wire [8:0] _T_405;
  wire [15:0] _GEN_48;
  wire [15:0] _T_406;
  wire [31:0] _GEN_49;
  wire [32:0] _T_407;
  wire [31:0] _T_408;
  wire [15:0] _T_410;
  wire [22:0] _GEN_50;
  wire [22:0] _T_411;
  wire [14:0] _T_412;
  wire  _T_416;
  wire [31:0] _GEN_51;
  wire [31:0] _T_417;
  wire [31:0] _T_418;
  wire [31:0] _T_419;
  wire [31:0] _T_420;
  wire [31:0] _T_421;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire  _T_424;
  wire  _T_425;
  wire [31:0] _T_426;
  wire [9:0] _T_429;
  wire [2:0] _T_430;
  wire [2:0] _T_431;
  wire [31:0] _GEN_53;
  wire [31:0] _T_432;
  wire [31:0] _T_433;
  wire  _T_434;
  wire  _T_436;
  wire [8:0] _GEN_54;
  wire [9:0] _T_437;
  wire [9:0] _T_438;
  wire [8:0] _T_439;
  wire  _GEN_8;
  wire [31:0] _GEN_9;
  wire [8:0] _GEN_10;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [7:0] Queue_2_io_enq_bits_strb;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [7:0] Queue_2_io_deq_bits_strb;
  wire  Queue_2_io_deq_bits_last;
  wire  _T_445_valid;
  wire [63:0] _T_445_bits_data;
  wire [7:0] _T_445_bits_strb;
  wire  _T_445_bits_last;
  wire [7:0] _T_449;
  reg  _T_452;
  reg [31:0] _RAND_6;
  wire  _T_457;
  wire  _GEN_11;
  wire  _T_459;
  wire  _GEN_12;
  wire  _T_461;
  wire  _T_462;
  wire  _T_464;
  wire  _T_466;
  wire  _T_467;
  wire [7:0] _T_468;
  reg [8:0] _T_471;
  reg [31:0] _RAND_7;
  wire  _T_473;
  wire [8:0] _T_475;
  wire [8:0] _T_476;
  wire  _T_478;
  wire  _T_479;
  wire [8:0] _GEN_55;
  wire [9:0] _T_480;
  wire [9:0] _T_481;
  wire [8:0] _T_482;
  wire  _T_485;
  wire  _T_487;
  wire  _T_488;
  wire  _T_489;
  wire  _T_491;
  wire  _T_493;
  wire  _T_494;
  wire  _T_495;
  wire  _T_499;
  wire  _T_501;
  wire  _T_503;
  wire  _T_504;
  wire  _T_505;
  wire  _T_506;
  wire  _T_508;
  wire  _T_512;
  wire  _T_515;
  wire  _T_516;
  Queue_32 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst),
    .io_deq_bits_user(Queue_io_deq_bits_user)
  );
  Queue_32 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_enq_bits_user(Queue_1_io_enq_bits_user),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst),
    .io_deq_bits_user(Queue_1_io_deq_bits_user)
  );
  Queue_11 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_strb(Queue_2_io_enq_bits_strb),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_strb(Queue_2_io_deq_bits_strb),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  assign io_out_0_aw_valid = _T_462;
  assign io_out_0_aw_bits_id = _T_273_bits_id;
  assign io_out_0_aw_bits_addr = _T_433;
  assign io_out_0_aw_bits_len = _T_398;
  assign io_out_0_aw_bits_size = _T_273_bits_size;
  assign io_out_0_aw_bits_user = _T_468;
  assign io_out_0_w_valid = _T_495;
  assign io_out_0_w_bits_data = _T_445_bits_data;
  assign io_out_0_w_bits_strb = _T_445_bits_strb;
  assign io_out_0_w_bits_last = _T_478;
  assign io_out_0_b_ready = _T_516;
  assign io_out_0_ar_valid = _T_95_valid;
  assign io_out_0_ar_bits_id = _T_95_bits_id;
  assign io_out_0_ar_bits_addr = _T_261;
  assign io_out_0_ar_bits_len = _T_226;
  assign io_out_0_ar_bits_size = _T_95_bits_size;
  assign io_out_0_ar_bits_user = _T_449;
  assign io_out_0_r_ready = io_in_0_r_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_ar_valid;
  assign Queue_io_enq_bits_id = io_in_0_ar_bits_id;
  assign Queue_io_enq_bits_addr = io_in_0_ar_bits_addr;
  assign Queue_io_enq_bits_len = io_in_0_ar_bits_len;
  assign Queue_io_enq_bits_size = io_in_0_ar_bits_size;
  assign Queue_io_enq_bits_burst = io_in_0_ar_bits_burst;
  assign Queue_io_enq_bits_user = io_in_0_ar_bits_user;
  assign Queue_io_deq_ready = _T_253;
  assign _T_95_valid = Queue_io_deq_valid;
  assign _T_95_bits_id = Queue_io_deq_bits_id;
  assign _T_95_bits_addr = Queue_io_deq_bits_addr;
  assign _T_95_bits_len = Queue_io_deq_bits_len;
  assign _T_95_bits_size = Queue_io_deq_bits_size;
  assign _T_95_bits_burst = Queue_io_deq_bits_burst;
  assign _T_95_bits_user = Queue_io_deq_bits_user;
  assign _T_110 = _T_105 ? _T_109 : _T_95_bits_len;
  assign _T_111 = _T_105 ? _T_107 : _T_95_bits_addr;
  assign _T_113 = _T_111[31:3];
  assign _T_114 = _T_113[7:0];
  assign _T_116 = _T_111 ^ 32'hc000000;
  assign _T_117 = {1'b0,$signed(_T_116)};
  assign _T_119 = $signed(_T_117) & $signed(33'shfc000000);
  assign _T_120 = $signed(_T_119);
  assign _T_122 = $signed(_T_120) == $signed(33'sh0);
  assign _T_124 = _T_111 ^ 32'h2000000;
  assign _T_125 = {1'b0,$signed(_T_124)};
  assign _T_127 = $signed(_T_125) & $signed(33'shffff0000);
  assign _T_128 = $signed(_T_127);
  assign _T_130 = $signed(_T_128) == $signed(33'sh0);
  assign _T_133 = {1'b0,$signed(_T_111)};
  assign _T_135 = $signed(_T_133) & $signed(33'shffffd000);
  assign _T_136 = $signed(_T_135);
  assign _T_138 = $signed(_T_136) == $signed(33'sh0);
  assign _T_140 = _T_111 ^ 32'h10000;
  assign _T_141 = {1'b0,$signed(_T_140)};
  assign _T_143 = $signed(_T_141) & $signed(33'shffff0000);
  assign _T_144 = $signed(_T_143);
  assign _T_146 = $signed(_T_144) == $signed(33'sh0);
  assign _T_148 = _T_111 ^ 32'h80000000;
  assign _T_149 = {1'b0,$signed(_T_148)};
  assign _T_151 = $signed(_T_149) & $signed(33'shffffc000);
  assign _T_152 = $signed(_T_151);
  assign _T_154 = $signed(_T_152) == $signed(33'sh0);
  assign _T_156 = _T_111 ^ 32'h60000000;
  assign _T_157 = {1'b0,$signed(_T_156)};
  assign _T_159 = $signed(_T_157) & $signed(33'she0000000);
  assign _T_160 = $signed(_T_159);
  assign _T_162 = $signed(_T_160) == $signed(33'sh0);
  assign _T_163 = _T_122 | _T_130;
  assign _T_164 = _T_163 | _T_138;
  assign _T_165 = _T_164 | _T_146;
  assign _T_166 = _T_165 | _T_154;
  assign _T_167 = _T_166 | _T_162;
  assign _T_170 = _T_111 ^ 32'h1000;
  assign _T_171 = {1'b0,$signed(_T_170)};
  assign _T_173 = $signed(_T_171) & $signed(33'shffffd000);
  assign _T_174 = $signed(_T_173);
  assign _T_176 = $signed(_T_174) == $signed(33'sh0);
  assign _T_180 = _T_167 ? 3'h7 : 3'h0;
  assign _T_182 = _T_176 ? 8'hff : 8'h0;
  assign _GEN_16 = {{5'd0}, _T_180};
  assign _T_183 = _GEN_16 | _T_182;
  assign _T_186 = _T_110[7:1];
  assign _GEN_17 = {{1'd0}, _T_186};
  assign _T_187 = _T_110 | _GEN_17;
  assign _T_188 = _T_187[7:2];
  assign _GEN_18 = {{2'd0}, _T_188};
  assign _T_189 = _T_187 | _GEN_18;
  assign _T_190 = _T_189[7:4];
  assign _GEN_19 = {{4'd0}, _T_190};
  assign _T_191 = _T_189 | _GEN_19;
  assign _T_193 = _T_191[7:1];
  assign _T_194 = ~ _T_110;
  assign _GEN_20 = {{1'd0}, _T_194};
  assign _T_195 = _GEN_20 << 1;
  assign _T_196 = _T_195[7:0];
  assign _T_197 = _T_194 | _T_196;
  assign _GEN_21 = {{2'd0}, _T_197};
  assign _T_198 = _GEN_21 << 2;
  assign _T_199 = _T_198[7:0];
  assign _T_200 = _T_197 | _T_199;
  assign _GEN_22 = {{4'd0}, _T_200};
  assign _T_201 = _GEN_22 << 4;
  assign _T_202 = _T_201[7:0];
  assign _T_203 = _T_200 | _T_202;
  assign _T_205 = ~ _T_203;
  assign _GEN_23 = {{1'd0}, _T_193};
  assign _T_206 = _GEN_23 | _T_205;
  assign _GEN_24 = {{1'd0}, _T_114};
  assign _T_207 = _GEN_24 << 1;
  assign _T_208 = _T_207[7:0];
  assign _T_209 = _T_114 | _T_208;
  assign _GEN_25 = {{2'd0}, _T_209};
  assign _T_210 = _GEN_25 << 2;
  assign _T_211 = _T_210[7:0];
  assign _T_212 = _T_209 | _T_211;
  assign _GEN_26 = {{4'd0}, _T_212};
  assign _T_213 = _GEN_26 << 4;
  assign _T_214 = _T_213[7:0];
  assign _T_215 = _T_212 | _T_214;
  assign _T_217 = ~ _T_215;
  assign _T_218 = _T_206 & _T_217;
  assign _T_219 = _T_218 & _T_183;
  assign _T_221 = _T_95_bits_burst == 2'h0;
  assign _T_223 = _T_95_bits_size != 3'h3;
  assign _T_224 = _T_221 | _T_223;
  assign _T_226 = _T_224 ? 8'h0 : _T_219;
  assign _GEN_27 = {{1'd0}, _T_226};
  assign _T_227 = _GEN_27 << 1;
  assign _T_229 = _T_227 | 9'h1;
  assign _T_231 = {1'h0,_T_226};
  assign _T_232 = ~ _T_231;
  assign _T_233 = _T_229 & _T_232;
  assign _GEN_28 = {{7'd0}, _T_233};
  assign _T_234 = _GEN_28 << _T_95_bits_size;
  assign _GEN_29 = {{16'd0}, _T_234};
  assign _T_235 = _T_111 + _GEN_29;
  assign _T_236 = _T_235[31:0];
  assign _T_238 = {_T_95_bits_len,8'hff};
  assign _GEN_30 = {{7'd0}, _T_238};
  assign _T_239 = _GEN_30 << _T_95_bits_size;
  assign _T_240 = _T_239[22:8];
  assign _T_244 = _T_95_bits_burst == 2'h2;
  assign _GEN_31 = {{17'd0}, _T_240};
  assign _T_245 = _T_236 & _GEN_31;
  assign _T_246 = ~ _T_95_bits_addr;
  assign _T_247 = _T_246 | _GEN_31;
  assign _T_248 = ~ _T_247;
  assign _T_249 = _T_245 | _T_248;
  assign _GEN_1 = _T_244 ? _T_249 : _T_236;
  assign _GEN_2 = _T_221 ? _T_95_bits_addr : _GEN_1;
  assign _T_252 = _T_226 == _T_110;
  assign _T_253 = io_out_0_ar_ready & _T_252;
  assign _T_254 = ~ _T_111;
  assign _T_257 = 10'h7 << _T_95_bits_size;
  assign _T_258 = _T_257[2:0];
  assign _T_259 = ~ _T_258;
  assign _GEN_33 = {{29'd0}, _T_259};
  assign _T_260 = _T_254 | _GEN_33;
  assign _T_261 = ~ _T_260;
  assign _T_262 = io_out_0_ar_ready & _T_95_valid;
  assign _T_264 = _T_252 == 1'h0;
  assign _GEN_34 = {{1'd0}, _T_110};
  assign _T_265 = _GEN_34 - _T_233;
  assign _T_266 = $unsigned(_T_265);
  assign _T_267 = _T_266[8:0];
  assign _GEN_3 = _T_262 ? _T_264 : _T_105;
  assign _GEN_4 = _T_262 ? _GEN_2 : _T_107;
  assign _GEN_5 = _T_262 ? _T_267 : {{1'd0}, _T_109};
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_in_0_aw_valid;
  assign Queue_1_io_enq_bits_id = io_in_0_aw_bits_id;
  assign Queue_1_io_enq_bits_addr = io_in_0_aw_bits_addr;
  assign Queue_1_io_enq_bits_len = io_in_0_aw_bits_len;
  assign Queue_1_io_enq_bits_size = io_in_0_aw_bits_size;
  assign Queue_1_io_enq_bits_burst = io_in_0_aw_bits_burst;
  assign Queue_1_io_enq_bits_user = io_in_0_aw_bits_user;
  assign Queue_1_io_deq_ready = _T_425;
  assign _T_273_valid = Queue_1_io_deq_valid;
  assign _T_273_bits_id = Queue_1_io_deq_bits_id;
  assign _T_273_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_273_bits_len = Queue_1_io_deq_bits_len;
  assign _T_273_bits_size = Queue_1_io_deq_bits_size;
  assign _T_273_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_273_bits_user = Queue_1_io_deq_bits_user;
  assign _T_288 = _T_283 ? _T_287 : _T_273_bits_len;
  assign _T_289 = _T_283 ? _T_285 : _T_273_bits_addr;
  assign _T_291 = _T_289[31:3];
  assign _T_292 = _T_291[7:0];
  assign _T_294 = _T_289 ^ 32'h60000000;
  assign _T_295 = {1'b0,$signed(_T_294)};
  assign _T_297 = $signed(_T_295) & $signed(33'she0000000);
  assign _T_298 = $signed(_T_297);
  assign _T_300 = $signed(_T_298) == $signed(33'sh0);
  assign _T_303 = _T_289 ^ 32'hc000000;
  assign _T_304 = {1'b0,$signed(_T_303)};
  assign _T_306 = $signed(_T_304) & $signed(33'shfc000000);
  assign _T_307 = $signed(_T_306);
  assign _T_309 = $signed(_T_307) == $signed(33'sh0);
  assign _T_311 = _T_289 ^ 32'h2000000;
  assign _T_312 = {1'b0,$signed(_T_311)};
  assign _T_314 = $signed(_T_312) & $signed(33'shffff0000);
  assign _T_315 = $signed(_T_314);
  assign _T_317 = $signed(_T_315) == $signed(33'sh0);
  assign _T_320 = {1'b0,$signed(_T_289)};
  assign _T_322 = $signed(_T_320) & $signed(33'shffffd000);
  assign _T_323 = $signed(_T_322);
  assign _T_325 = $signed(_T_323) == $signed(33'sh0);
  assign _T_327 = _T_289 ^ 32'h80000000;
  assign _T_328 = {1'b0,$signed(_T_327)};
  assign _T_330 = $signed(_T_328) & $signed(33'shffffc000);
  assign _T_331 = $signed(_T_330);
  assign _T_333 = $signed(_T_331) == $signed(33'sh0);
  assign _T_334 = _T_309 | _T_317;
  assign _T_335 = _T_334 | _T_325;
  assign _T_336 = _T_335 | _T_333;
  assign _T_339 = _T_289 ^ 32'h1000;
  assign _T_340 = {1'b0,$signed(_T_339)};
  assign _T_342 = $signed(_T_340) & $signed(33'shffffd000);
  assign _T_343 = $signed(_T_342);
  assign _T_345 = $signed(_T_343) == $signed(33'sh0);
  assign _T_349 = _T_300 ? 5'h1f : 5'h0;
  assign _T_351 = _T_336 ? 3'h7 : 3'h0;
  assign _T_353 = _T_345 ? 8'hff : 8'h0;
  assign _GEN_35 = {{2'd0}, _T_351};
  assign _T_354 = _T_349 | _GEN_35;
  assign _GEN_36 = {{3'd0}, _T_354};
  assign _T_355 = _GEN_36 | _T_353;
  assign _T_358 = _T_288[7:1];
  assign _GEN_37 = {{1'd0}, _T_358};
  assign _T_359 = _T_288 | _GEN_37;
  assign _T_360 = _T_359[7:2];
  assign _GEN_38 = {{2'd0}, _T_360};
  assign _T_361 = _T_359 | _GEN_38;
  assign _T_362 = _T_361[7:4];
  assign _GEN_39 = {{4'd0}, _T_362};
  assign _T_363 = _T_361 | _GEN_39;
  assign _T_365 = _T_363[7:1];
  assign _T_366 = ~ _T_288;
  assign _GEN_40 = {{1'd0}, _T_366};
  assign _T_367 = _GEN_40 << 1;
  assign _T_368 = _T_367[7:0];
  assign _T_369 = _T_366 | _T_368;
  assign _GEN_41 = {{2'd0}, _T_369};
  assign _T_370 = _GEN_41 << 2;
  assign _T_371 = _T_370[7:0];
  assign _T_372 = _T_369 | _T_371;
  assign _GEN_42 = {{4'd0}, _T_372};
  assign _T_373 = _GEN_42 << 4;
  assign _T_374 = _T_373[7:0];
  assign _T_375 = _T_372 | _T_374;
  assign _T_377 = ~ _T_375;
  assign _GEN_43 = {{1'd0}, _T_365};
  assign _T_378 = _GEN_43 | _T_377;
  assign _GEN_44 = {{1'd0}, _T_292};
  assign _T_379 = _GEN_44 << 1;
  assign _T_380 = _T_379[7:0];
  assign _T_381 = _T_292 | _T_380;
  assign _GEN_45 = {{2'd0}, _T_381};
  assign _T_382 = _GEN_45 << 2;
  assign _T_383 = _T_382[7:0];
  assign _T_384 = _T_381 | _T_383;
  assign _GEN_46 = {{4'd0}, _T_384};
  assign _T_385 = _GEN_46 << 4;
  assign _T_386 = _T_385[7:0];
  assign _T_387 = _T_384 | _T_386;
  assign _T_389 = ~ _T_387;
  assign _T_390 = _T_378 & _T_389;
  assign _T_391 = _T_390 & _T_355;
  assign _T_393 = _T_273_bits_burst == 2'h0;
  assign _T_395 = _T_273_bits_size != 3'h3;
  assign _T_396 = _T_393 | _T_395;
  assign _T_398 = _T_396 ? 8'h0 : _T_391;
  assign _GEN_47 = {{1'd0}, _T_398};
  assign _T_399 = _GEN_47 << 1;
  assign _T_401 = _T_399 | 9'h1;
  assign _T_403 = {1'h0,_T_398};
  assign _T_404 = ~ _T_403;
  assign _T_405 = _T_401 & _T_404;
  assign _GEN_48 = {{7'd0}, _T_405};
  assign _T_406 = _GEN_48 << _T_273_bits_size;
  assign _GEN_49 = {{16'd0}, _T_406};
  assign _T_407 = _T_289 + _GEN_49;
  assign _T_408 = _T_407[31:0];
  assign _T_410 = {_T_273_bits_len,8'hff};
  assign _GEN_50 = {{7'd0}, _T_410};
  assign _T_411 = _GEN_50 << _T_273_bits_size;
  assign _T_412 = _T_411[22:8];
  assign _T_416 = _T_273_bits_burst == 2'h2;
  assign _GEN_51 = {{17'd0}, _T_412};
  assign _T_417 = _T_408 & _GEN_51;
  assign _T_418 = ~ _T_273_bits_addr;
  assign _T_419 = _T_418 | _GEN_51;
  assign _T_420 = ~ _T_419;
  assign _T_421 = _T_417 | _T_420;
  assign _GEN_6 = _T_416 ? _T_421 : _T_408;
  assign _GEN_7 = _T_393 ? _T_273_bits_addr : _GEN_6;
  assign _T_424 = _T_398 == _T_288;
  assign _T_425 = _T_464 & _T_424;
  assign _T_426 = ~ _T_289;
  assign _T_429 = 10'h7 << _T_273_bits_size;
  assign _T_430 = _T_429[2:0];
  assign _T_431 = ~ _T_430;
  assign _GEN_53 = {{29'd0}, _T_431};
  assign _T_432 = _T_426 | _GEN_53;
  assign _T_433 = ~ _T_432;
  assign _T_434 = _T_464 & _T_273_valid;
  assign _T_436 = _T_424 == 1'h0;
  assign _GEN_54 = {{1'd0}, _T_288};
  assign _T_437 = _GEN_54 - _T_405;
  assign _T_438 = $unsigned(_T_437);
  assign _T_439 = _T_438[8:0];
  assign _GEN_8 = _T_434 ? _T_436 : _T_283;
  assign _GEN_9 = _T_434 ? _GEN_7 : _T_285;
  assign _GEN_10 = _T_434 ? _T_439 : {{1'd0}, _T_287};
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = io_in_0_w_valid;
  assign Queue_2_io_enq_bits_data = io_in_0_w_bits_data;
  assign Queue_2_io_enq_bits_strb = io_in_0_w_bits_strb;
  assign Queue_2_io_enq_bits_last = io_in_0_w_bits_last;
  assign Queue_2_io_deq_ready = _T_499;
  assign _T_445_valid = Queue_2_io_deq_valid;
  assign _T_445_bits_data = Queue_2_io_deq_bits_data;
  assign _T_445_bits_strb = Queue_2_io_deq_bits_strb;
  assign _T_445_bits_last = Queue_2_io_deq_bits_last;
  assign _T_449 = {_T_95_bits_user,_T_252};
  assign _T_457 = _T_467 & _T_473;
  assign _GEN_11 = _T_457 ? 1'h1 : _T_452;
  assign _T_459 = io_out_0_aw_ready & io_out_0_aw_valid;
  assign _GEN_12 = _T_459 ? 1'h0 : _GEN_11;
  assign _T_461 = _T_473 | _T_452;
  assign _T_462 = _T_273_valid & _T_461;
  assign _T_464 = io_out_0_aw_ready & _T_461;
  assign _T_466 = _T_452 == 1'h0;
  assign _T_467 = _T_273_valid & _T_466;
  assign _T_468 = {_T_273_bits_user,_T_424};
  assign _T_473 = _T_471 == 9'h0;
  assign _T_475 = _T_467 ? _T_405 : 9'h0;
  assign _T_476 = _T_473 ? _T_475 : _T_471;
  assign _T_478 = _T_476 == 9'h1;
  assign _T_479 = io_out_0_w_ready & io_out_0_w_valid;
  assign _GEN_55 = {{8'd0}, _T_479};
  assign _T_480 = _T_476 - _GEN_55;
  assign _T_481 = $unsigned(_T_480);
  assign _T_482 = _T_481[8:0];
  assign _T_485 = _T_479 == 1'h0;
  assign _T_487 = _T_476 != 9'h0;
  assign _T_488 = _T_485 | _T_487;
  assign _T_489 = _T_488 | reset;
  assign _T_491 = _T_489 == 1'h0;
  assign _T_493 = _T_473 == 1'h0;
  assign _T_494 = _T_493 | _T_467;
  assign _T_495 = _T_445_valid & _T_494;
  assign _T_499 = io_out_0_w_ready & _T_494;
  assign _T_501 = io_out_0_w_valid == 1'h0;
  assign _T_503 = _T_445_bits_last == 1'h0;
  assign _T_504 = _T_501 | _T_503;
  assign _T_505 = _T_504 | _T_478;
  assign _T_506 = _T_505 | reset;
  assign _T_508 = _T_506 == 1'h0;
  assign _T_512 = io_out_0_b_bits_user[0];
  assign _T_515 = _T_512 == 1'h0;
  assign _T_516 = io_in_0_b_ready | _T_515;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_105 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_107 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_109 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_283 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_285 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_287 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_452 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_471 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_105 <= 1'h0;
    end else begin
      if (_T_262) begin
        _T_105 <= _T_264;
      end
    end
    if (_T_262) begin
      if (_T_221) begin
        _T_107 <= _T_95_bits_addr;
      end else begin
        if (_T_244) begin
          _T_107 <= _T_249;
        end else begin
          _T_107 <= _T_236;
        end
      end
    end
    _T_109 <= _GEN_5[7:0];
    if (reset) begin
      _T_283 <= 1'h0;
    end else begin
      if (_T_434) begin
        _T_283 <= _T_436;
      end
    end
    if (_T_434) begin
      if (_T_393) begin
        _T_285 <= _T_273_bits_addr;
      end else begin
        if (_T_416) begin
          _T_285 <= _T_421;
        end else begin
          _T_285 <= _T_408;
        end
      end
    end
    _T_287 <= _GEN_10[7:0];
    if (reset) begin
      _T_452 <= 1'h0;
    end else begin
      if (_T_459) begin
        _T_452 <= 1'h0;
      end else begin
        if (_T_457) begin
          _T_452 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_471 <= 9'h0;
    end else begin
      _T_471 <= _T_482;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_491) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:172 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_491) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_508) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:181 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_508) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_35(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
  reg [7:0] ram [0:3];
  reg [31:0] _RAND_0;
  wire [7:0] ram__T_43_data;
  wire [1:0] ram__T_43_addr;
  wire [7:0] ram__T_29_data;
  wire [1:0] ram__T_29_addr;
  wire  ram__T_29_mask;
  wire  ram__T_29_en;
  reg [1:0] value;
  reg [31:0] _RAND_1;
  reg [1:0] value_1;
  reg [31:0] _RAND_2;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [2:0] _T_32;
  wire [1:0] _T_33;
  wire [1:0] _GEN_4;
  wire [2:0] _T_36;
  wire [1:0] _T_37;
  wire [1:0] _GEN_5;
  wire  _T_38;
  wire  _GEN_6;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits = ram__T_43_data;
  assign ram__T_43_addr = value_1;
  assign ram__T_43_data = ram[ram__T_43_addr];
  assign ram__T_29_data = io_enq_bits;
  assign ram__T_29_addr = value;
  assign ram__T_29_mask = _T_25;
  assign ram__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 2'h1;
  assign _T_33 = _T_32[1:0];
  assign _GEN_4 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 2'h1;
  assign _T_37 = _T_36[1:0];
  assign _GEN_5 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_6 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  value = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  value_1 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram__T_29_en & ram__T_29_mask) begin
      ram[ram__T_29_addr] <= ram__T_29_data;
    end
    if (reset) begin
      value <= 2'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module AXI4UserYanker_1(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input         io_in_0_aw_bits_id,
  input  [31:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [7:0]  io_in_0_aw_bits_user,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output [7:0]  io_in_0_b_bits_user,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input         io_in_0_ar_bits_id,
  input  [31:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [7:0]  io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output        io_out_0_aw_bits_id,
  output [31:0] io_out_0_aw_bits_addr,
  output [7:0]  io_out_0_aw_bits_len,
  output [2:0]  io_out_0_aw_bits_size,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input         io_out_0_b_bits_id,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output        io_out_0_ar_bits_id,
  output [31:0] io_out_0_ar_bits_addr,
  output [7:0]  io_out_0_ar_bits_len,
  output [2:0]  io_out_0_ar_bits_size,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input         io_out_0_r_bits_id,
  input         io_out_0_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [7:0] Queue_io_enq_bits;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [7:0] Queue_io_deq_bits;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [7:0] Queue_1_io_enq_bits;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [7:0] Queue_1_io_deq_bits;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [7:0] Queue_2_io_enq_bits;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [7:0] Queue_2_io_deq_bits;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [7:0] Queue_3_io_enq_bits;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [7:0] Queue_3_io_deq_bits;
  wire  _T_96_0;
  wire  _T_96_1;
  wire  _GEN_8;
  wire  _T_102;
  wire  _T_103;
  wire  _T_106_0;
  wire  _T_106_1;
  wire  _T_121;
  wire  _GEN_9;
  wire  _T_122;
  wire  _T_123;
  wire  _T_125;
  wire [1:0] _T_128;
  wire  _T_130;
  wire  _T_131;
  wire [1:0] _T_134;
  wire  _T_136;
  wire  _T_137;
  wire  _T_138;
  wire  _T_139;
  wire  _T_140;
  wire  _T_141;
  wire  _T_142;
  wire  _T_144;
  wire  _T_145;
  wire  _T_147;
  wire  _T_150_0;
  wire  _T_150_1;
  wire  _GEN_11;
  wire  _T_156;
  wire  _T_157;
  wire  _T_160_0;
  wire  _T_160_1;
  wire [7:0] _T_168_0;
  wire [7:0] _T_168_1;
  wire  _T_175;
  wire  _GEN_12;
  wire  _T_176;
  wire  _T_177;
  wire  _T_179;
  wire [7:0] _GEN_13;
  wire [1:0] _T_182;
  wire  _T_184;
  wire  _T_185;
  wire [1:0] _T_188;
  wire  _T_190;
  wire  _T_191;
  wire  _T_192;
  wire  _T_193;
  wire  _T_194;
  wire  _T_195;
  wire  _T_197;
  wire  _T_199;
  Queue_35 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits(Queue_io_enq_bits),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits(Queue_io_deq_bits)
  );
  Queue_35 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits(Queue_1_io_enq_bits),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits(Queue_1_io_deq_bits)
  );
  Queue_35 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits(Queue_2_io_enq_bits),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits(Queue_2_io_deq_bits)
  );
  Queue_35 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits(Queue_3_io_enq_bits),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits(Queue_3_io_deq_bits)
  );
  assign io_in_0_aw_ready = _T_156;
  assign io_in_0_w_ready = io_out_0_w_ready;
  assign io_in_0_b_bits_user = _GEN_13;
  assign io_in_0_ar_ready = _T_102;
  assign io_out_0_aw_valid = _T_157;
  assign io_out_0_aw_bits_id = io_in_0_aw_bits_id;
  assign io_out_0_aw_bits_addr = io_in_0_aw_bits_addr;
  assign io_out_0_aw_bits_len = io_in_0_aw_bits_len;
  assign io_out_0_aw_bits_size = io_in_0_aw_bits_size;
  assign io_out_0_w_valid = io_in_0_w_valid;
  assign io_out_0_w_bits_data = io_in_0_w_bits_data;
  assign io_out_0_w_bits_strb = io_in_0_w_bits_strb;
  assign io_out_0_w_bits_last = io_in_0_w_bits_last;
  assign io_out_0_b_ready = io_in_0_b_ready;
  assign io_out_0_ar_valid = _T_103;
  assign io_out_0_ar_bits_id = io_in_0_ar_bits_id;
  assign io_out_0_ar_bits_addr = io_in_0_ar_bits_addr;
  assign io_out_0_ar_bits_len = io_in_0_ar_bits_len;
  assign io_out_0_ar_bits_size = io_in_0_ar_bits_size;
  assign io_out_0_r_ready = io_in_0_r_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_142;
  assign Queue_io_enq_bits = io_in_0_ar_bits_user;
  assign Queue_io_deq_ready = _T_140;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_147;
  assign Queue_1_io_enq_bits = io_in_0_ar_bits_user;
  assign Queue_1_io_deq_ready = _T_145;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = _T_195;
  assign Queue_2_io_enq_bits = io_in_0_aw_bits_user;
  assign Queue_2_io_deq_ready = _T_193;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = _T_199;
  assign Queue_3_io_enq_bits = io_in_0_aw_bits_user;
  assign Queue_3_io_deq_ready = _T_197;
  assign _T_96_0 = Queue_io_enq_ready;
  assign _T_96_1 = Queue_1_io_enq_ready;
  assign _GEN_8 = io_in_0_ar_bits_id ? _T_96_1 : _T_96_0;
  assign _T_102 = io_out_0_ar_ready & _GEN_8;
  assign _T_103 = io_in_0_ar_valid & _GEN_8;
  assign _T_106_0 = Queue_io_deq_valid;
  assign _T_106_1 = Queue_1_io_deq_valid;
  assign _T_121 = io_out_0_r_valid == 1'h0;
  assign _GEN_9 = io_out_0_r_bits_id ? _T_106_1 : _T_106_0;
  assign _T_122 = _T_121 | _GEN_9;
  assign _T_123 = _T_122 | reset;
  assign _T_125 = _T_123 == 1'h0;
  assign _T_128 = 2'h1 << io_in_0_ar_bits_id;
  assign _T_130 = _T_128[0];
  assign _T_131 = _T_128[1];
  assign _T_134 = 2'h1 << io_out_0_r_bits_id;
  assign _T_136 = _T_134[0];
  assign _T_137 = _T_134[1];
  assign _T_138 = io_out_0_r_valid & io_in_0_r_ready;
  assign _T_139 = _T_138 & _T_136;
  assign _T_140 = _T_139 & io_out_0_r_bits_last;
  assign _T_141 = io_in_0_ar_valid & io_out_0_ar_ready;
  assign _T_142 = _T_141 & _T_130;
  assign _T_144 = _T_138 & _T_137;
  assign _T_145 = _T_144 & io_out_0_r_bits_last;
  assign _T_147 = _T_141 & _T_131;
  assign _T_150_0 = Queue_2_io_enq_ready;
  assign _T_150_1 = Queue_3_io_enq_ready;
  assign _GEN_11 = io_in_0_aw_bits_id ? _T_150_1 : _T_150_0;
  assign _T_156 = io_out_0_aw_ready & _GEN_11;
  assign _T_157 = io_in_0_aw_valid & _GEN_11;
  assign _T_160_0 = Queue_2_io_deq_valid;
  assign _T_160_1 = Queue_3_io_deq_valid;
  assign _T_168_0 = Queue_2_io_deq_bits;
  assign _T_168_1 = Queue_3_io_deq_bits;
  assign _T_175 = io_out_0_b_valid == 1'h0;
  assign _GEN_12 = io_out_0_b_bits_id ? _T_160_1 : _T_160_0;
  assign _T_176 = _T_175 | _GEN_12;
  assign _T_177 = _T_176 | reset;
  assign _T_179 = _T_177 == 1'h0;
  assign _GEN_13 = io_out_0_b_bits_id ? _T_168_1 : _T_168_0;
  assign _T_182 = 2'h1 << io_in_0_aw_bits_id;
  assign _T_184 = _T_182[0];
  assign _T_185 = _T_182[1];
  assign _T_188 = 2'h1 << io_out_0_b_bits_id;
  assign _T_190 = _T_188[0];
  assign _T_191 = _T_188[1];
  assign _T_192 = io_out_0_b_valid & io_in_0_b_ready;
  assign _T_193 = _T_192 & _T_190;
  assign _T_194 = io_in_0_aw_valid & io_out_0_aw_ready;
  assign _T_195 = _T_194 & _T_184;
  assign _T_197 = _T_192 & _T_191;
  assign _T_199 = _T_194 & _T_185;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_125) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:60 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_125) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_179) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UserYanker.scala:81 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_179) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_39(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_id,
  input   io_enq_bits_last,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_id,
  output  io_deq_bits_last
);
  reg  ram_id [0:0];
  reg [31:0] _RAND_0;
  wire  ram_id__T_35_data;
  wire  ram_id__T_35_addr;
  wire  ram_id__T_26_data;
  wire  ram_id__T_26_addr;
  wire  ram_id__T_26_mask;
  wire  ram_id__T_26_en;
  reg  ram_last [0:0];
  reg [31:0] _RAND_1;
  wire  ram_last__T_35_data;
  wire  ram_last__T_35_addr;
  wire  ram_last__T_26_data;
  wire  ram_last__T_26_addr;
  wire  ram_last__T_26_mask;
  wire  ram_last__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_2;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_7;
  wire  _T_31;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _GEN_10;
  wire  _GEN_13;
  wire  _GEN_14;
  wire  _GEN_15;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_8;
  assign io_deq_bits_id = _GEN_10;
  assign io_deq_bits_last = _GEN_13;
  assign ram_id__T_35_addr = 1'h0;
  assign ram_id__T_35_data = ram_id[ram_id__T_35_addr];
  assign ram_id__T_26_data = io_enq_bits_id;
  assign ram_id__T_26_addr = 1'h0;
  assign ram_id__T_26_mask = _GEN_15;
  assign ram_id__T_26_en = _GEN_15;
  assign ram_last__T_35_addr = 1'h0;
  assign ram_last__T_35_data = ram_last[ram_last__T_35_addr];
  assign ram_last__T_26_data = io_enq_bits_last;
  assign ram_last__T_26_addr = 1'h0;
  assign ram_last__T_26_mask = _GEN_15;
  assign ram_last__T_26_en = _GEN_15;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_15 != _GEN_14;
  assign _GEN_7 = _T_29 ? _GEN_15 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_8 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_9 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_10 = _T_18 ? io_enq_bits_id : ram_id__T_35_data;
  assign _GEN_13 = _T_18 ? io_enq_bits_last : ram_last__T_35_data;
  assign _GEN_14 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_15 = _T_18 ? _GEN_9 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_last[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  maybe_full = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_26_en & ram_id__T_26_mask) begin
      ram_id[ram_id__T_26_addr] <= ram_id__T_26_data;
    end
    if(ram_last__T_26_en & ram_last__T_26_mask) begin
      ram_last[ram_last__T_26_addr] <= ram_last__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module Queue_40(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits_id
);
  reg  ram_id [0:0];
  reg [31:0] _RAND_0;
  wire  ram_id__T_35_data;
  wire  ram_id__T_35_addr;
  wire  ram_id__T_26_data;
  wire  ram_id__T_26_addr;
  wire  ram_id__T_26_mask;
  wire  ram_id__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_1;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_5;
  wire  _T_31;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_10;
  wire  _GEN_11;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_6;
  assign io_deq_bits_id = _GEN_8;
  assign ram_id__T_35_addr = 1'h0;
  assign ram_id__T_35_data = ram_id[ram_id__T_35_addr];
  assign ram_id__T_26_data = io_enq_bits_id;
  assign ram_id__T_26_addr = 1'h0;
  assign ram_id__T_26_mask = _GEN_11;
  assign ram_id__T_26_en = _GEN_11;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_11 != _GEN_10;
  assign _GEN_5 = _T_29 ? _GEN_11 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_6 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_7 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_8 = _T_18 ? io_enq_bits_id : ram_id__T_35_data;
  assign _GEN_10 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_11 = _T_18 ? _GEN_7 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  maybe_full = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_26_en & ram_id__T_26_mask) begin
      ram_id[ram_id__T_26_addr] <= ram_id__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module AXI4ToTL(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input         io_in_0_aw_bits_id,
  input  [31:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output        io_in_0_b_bits_id,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input         io_in_0_ar_bits_id,
  input  [31:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output        io_in_0_r_bits_id,
  output        io_in_0_r_bits_last,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output [3:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [7:0]  io_out_0_a_bits_mask,
  output [63:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input  [3:0]  io_out_0_d_bits_source
);
  wire [15:0] _T_95;
  wire [22:0] _GEN_16;
  wire [22:0] _T_96;
  wire [14:0] _T_97;
  wire [15:0] _GEN_17;
  wire [15:0] _T_98;
  wire [15:0] _T_100;
  wire [15:0] _T_102;
  wire [15:0] _T_103;
  wire [15:0] _T_104;
  wire [7:0] _T_105;
  wire [7:0] _T_106;
  wire  _T_108;
  wire [7:0] _T_109;
  wire [3:0] _T_110;
  wire [3:0] _T_111;
  wire  _T_113;
  wire [3:0] _T_114;
  wire [1:0] _T_115;
  wire [1:0] _T_116;
  wire  _T_118;
  wire [1:0] _T_119;
  wire  _T_120;
  wire [1:0] _T_121;
  wire [2:0] _T_122;
  wire [3:0] _T_123;
  wire  _T_128;
  wire [31:0] _T_132;
  wire [32:0] _T_133;
  wire [32:0] _T_135;
  wire [32:0] _T_136;
  wire  _T_138;
  wire  _T_139;
  wire  _T_144;
  wire [31:0] _T_148;
  wire [32:0] _T_149;
  wire [32:0] _T_151;
  wire [32:0] _T_152;
  wire  _T_154;
  wire [31:0] _T_156;
  wire [32:0] _T_157;
  wire [32:0] _T_159;
  wire [32:0] _T_160;
  wire  _T_162;
  wire [32:0] _T_165;
  wire [32:0] _T_167;
  wire [32:0] _T_168;
  wire  _T_170;
  wire [31:0] _T_172;
  wire [32:0] _T_173;
  wire [32:0] _T_175;
  wire [32:0] _T_176;
  wire  _T_178;
  wire [31:0] _T_180;
  wire [32:0] _T_181;
  wire [32:0] _T_183;
  wire [32:0] _T_184;
  wire  _T_186;
  wire [31:0] _T_188;
  wire [32:0] _T_189;
  wire [32:0] _T_191;
  wire [32:0] _T_192;
  wire  _T_194;
  wire  _T_195;
  wire  _T_196;
  wire  _T_197;
  wire  _T_198;
  wire  _T_199;
  wire  _T_200;
  wire  _T_203;
  wire [2:0] _T_205;
  wire [13:0] _GEN_18;
  wire [13:0] _T_206;
  wire [31:0] _T_207;
  reg [2:0] _T_225_0;
  reg [31:0] _RAND_0;
  reg [2:0] _T_225_1;
  reg [31:0] _RAND_1;
  wire [2:0] _GEN_4;
  wire [1:0] _T_239;
  wire [2:0] _T_241;
  wire [3:0] _T_242;
  wire  _T_244;
  wire [29:0] _T_247;
  wire [14:0] _T_248;
  wire [14:0] _T_249;
  wire  _T_250;
  wire  _T_251;
  wire  _T_252;
  wire  _T_254;
  wire [1:0] _T_339;
  wire [3:0] _T_341;
  wire [2:0] _T_342;
  wire [2:0] _T_344;
  wire  _T_346;
  wire  _T_348;
  wire  _T_349;
  wire  _T_351;
  wire  _T_353;
  wire  _T_354;
  wire  _T_356;
  wire  _T_357;
  wire  _T_358;
  wire  _T_359;
  wire  _T_361;
  wire  _T_362;
  wire  _T_363;
  wire  _T_364;
  wire  _T_365;
  wire  _T_366;
  wire  _T_367;
  wire  _T_368;
  wire  _T_369;
  wire  _T_370;
  wire  _T_371;
  wire  _T_372;
  wire  _T_373;
  wire  _T_374;
  wire  _T_375;
  wire  _T_377;
  wire  _T_378;
  wire  _T_379;
  wire  _T_380;
  wire  _T_381;
  wire  _T_382;
  wire  _T_383;
  wire  _T_384;
  wire  _T_385;
  wire  _T_386;
  wire  _T_387;
  wire  _T_388;
  wire  _T_389;
  wire  _T_390;
  wire  _T_391;
  wire  _T_392;
  wire  _T_393;
  wire  _T_394;
  wire  _T_395;
  wire  _T_396;
  wire  _T_397;
  wire  _T_398;
  wire  _T_399;
  wire  _T_400;
  wire  _T_401;
  wire [1:0] _T_402;
  wire [1:0] _T_403;
  wire [3:0] _T_404;
  wire [1:0] _T_405;
  wire [1:0] _T_406;
  wire [3:0] _T_407;
  wire [7:0] _T_408;
  wire [1:0] _T_412;
  wire  _T_414;
  wire  _T_415;
  wire  _T_416;
  wire  _T_417;
  wire [3:0] _T_419;
  wire [2:0] _T_420;
  wire [2:0] _GEN_5;
  wire  _T_422;
  wire [3:0] _T_424;
  wire [2:0] _T_425;
  wire [2:0] _GEN_6;
  wire [15:0] _T_431;
  wire [22:0] _GEN_19;
  wire [22:0] _T_432;
  wire [14:0] _T_433;
  wire [15:0] _GEN_20;
  wire [15:0] _T_434;
  wire [15:0] _T_436;
  wire [15:0] _T_438;
  wire [15:0] _T_439;
  wire [15:0] _T_440;
  wire [7:0] _T_441;
  wire [7:0] _T_442;
  wire  _T_444;
  wire [7:0] _T_445;
  wire [3:0] _T_446;
  wire [3:0] _T_447;
  wire  _T_449;
  wire [3:0] _T_450;
  wire [1:0] _T_451;
  wire [1:0] _T_452;
  wire  _T_454;
  wire [1:0] _T_455;
  wire  _T_456;
  wire [1:0] _T_457;
  wire [2:0] _T_458;
  wire [3:0] _T_459;
  wire  _T_464;
  wire [31:0] _T_468;
  wire [32:0] _T_469;
  wire [32:0] _T_471;
  wire [32:0] _T_472;
  wire  _T_474;
  wire  _T_475;
  wire  _T_480;
  wire [31:0] _T_484;
  wire [32:0] _T_485;
  wire [32:0] _T_487;
  wire [32:0] _T_488;
  wire  _T_490;
  wire [31:0] _T_492;
  wire [32:0] _T_493;
  wire [32:0] _T_495;
  wire [32:0] _T_496;
  wire  _T_498;
  wire [32:0] _T_501;
  wire [32:0] _T_503;
  wire [32:0] _T_504;
  wire  _T_506;
  wire [31:0] _T_508;
  wire [32:0] _T_509;
  wire [32:0] _T_511;
  wire [32:0] _T_512;
  wire  _T_514;
  wire  _T_515;
  wire  _T_516;
  wire  _T_517;
  wire  _T_518;
  wire  _T_523;
  wire [31:0] _T_527;
  wire [32:0] _T_528;
  wire [32:0] _T_530;
  wire [32:0] _T_531;
  wire  _T_533;
  wire  _T_534;
  wire  _T_549;
  wire  _T_550;
  wire [2:0] _T_553;
  wire [13:0] _GEN_21;
  wire [13:0] _T_554;
  wire [31:0] _T_555;
  reg [2:0] _T_573_0;
  reg [31:0] _RAND_2;
  reg [2:0] _T_573_1;
  reg [31:0] _RAND_3;
  wire [2:0] _GEN_7;
  wire [1:0] _T_587;
  wire [2:0] _T_589;
  wire [3:0] _T_590;
  wire  _T_592;
  wire [29:0] _T_595;
  wire [14:0] _T_596;
  wire [14:0] _T_597;
  wire  _T_598;
  wire  _T_599;
  wire  _T_600;
  wire  _T_602;
  wire  _T_606;
  wire  _T_607;
  wire  _T_609;
  wire  _T_610;
  wire  _T_611;
  wire  _T_613;
  wire  _T_614;
  wire  _T_615;
  wire  _T_616;
  wire  _T_617;
  wire [1:0] _T_716;
  wire  _T_718;
  wire  _T_719;
  wire  _T_720;
  wire  _T_721;
  wire [3:0] _T_723;
  wire [2:0] _T_724;
  wire [2:0] _GEN_8;
  wire  _T_726;
  wire [3:0] _T_728;
  wire [2:0] _T_729;
  wire [2:0] _GEN_9;
  reg [7:0] _T_733;
  reg [31:0] _RAND_4;
  wire  _T_735;
  wire  _T_736;
  wire [1:0] _T_737;
  wire  _T_739;
  wire  _T_740;
  wire  _T_742;
  reg [1:0] _T_746;
  reg [31:0] _RAND_5;
  wire [1:0] _T_747;
  wire [1:0] _T_748;
  wire [3:0] _T_749;
  wire [2:0] _T_750;
  wire [3:0] _GEN_22;
  wire [3:0] _T_751;
  wire [2:0] _T_753;
  wire [3:0] _GEN_23;
  wire [3:0] _T_754;
  wire [3:0] _GEN_24;
  wire [3:0] _T_755;
  wire [1:0] _T_756;
  wire [1:0] _T_757;
  wire [1:0] _T_758;
  wire [1:0] _T_759;
  wire  _T_761;
  wire  _T_762;
  wire [1:0] _T_763;
  wire [2:0] _GEN_25;
  wire [2:0] _T_764;
  wire [1:0] _T_765;
  wire [1:0] _T_766;
  wire [1:0] _GEN_10;
  wire  _T_769;
  wire  _T_770;
  wire  _T_778;
  wire  _T_779;
  wire  _T_789;
  wire  _T_793;
  wire  _T_798;
  wire  _T_799;
  wire  _T_801;
  wire  _T_803;
  wire  _T_804;
  wire  _T_806;
  wire  _T_808;
  wire  _T_809;
  wire  _T_811;
  wire [7:0] _T_815;
  wire  _T_817;
  wire [7:0] _GEN_26;
  wire [8:0] _T_818;
  wire [8:0] _T_819;
  wire [7:0] _T_820;
  wire [7:0] _T_821;
  reg  _T_839_0;
  reg [31:0] _RAND_6;
  reg  _T_839_1;
  reg [31:0] _RAND_7;
  wire  _T_850_0;
  wire  _T_850_1;
  wire  _T_858_0;
  wire  _T_858_1;
  wire  _T_866;
  wire  _T_867;
  wire  _T_871;
  wire  _T_873;
  wire  _T_874;
  wire  _T_877;
  wire [39:0] _T_879;
  wire [103:0] _T_880;
  wire [7:0] _T_881;
  wire [13:0] _T_883;
  wire [117:0] _T_884;
  wire [117:0] _T_886;
  wire [39:0] _T_887;
  wire [103:0] _T_888;
  wire [7:0] _T_889;
  wire [13:0] _T_891;
  wire [117:0] _T_892;
  wire [117:0] _T_894;
  wire [117:0] _T_895;
  wire [63:0] _T_900;
  wire [7:0] _T_901;
  wire [31:0] _T_902;
  wire [3:0] _T_903;
  wire [3:0] _T_904;
  wire [2:0] _T_905;
  wire [2:0] _T_906;
  wire  _T_907_ready;
  wire  _T_911_ready;
  wire  _T_918;
  wire  _T_919;
  wire [26:0] _T_922;
  wire [11:0] _T_923;
  wire [11:0] _T_924;
  wire [8:0] _T_925;
  wire [8:0] _T_928;
  reg [8:0] _T_931;
  reg [31:0] _RAND_8;
  wire [9:0] _T_933;
  wire [9:0] _T_934;
  wire [8:0] _T_935;
  wire  _T_937;
  wire  _T_939;
  wire  _T_941;
  wire  _T_942;
  wire [8:0] _T_946;
  wire [8:0] _GEN_11;
  wire  _T_947;
  wire  _T_948;
  wire  _T_950;
  wire  _T_951;
  wire  _T_952;
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire  Queue_io_enq_bits_id;
  wire  Queue_io_enq_bits_last;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire  Queue_io_deq_bits_id;
  wire  Queue_io_deq_bits_last;
  wire  _T_958_valid;
  wire  _T_958_bits_id;
  wire  _T_958_bits_last;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire  Queue_1_io_enq_bits_id;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire  Queue_1_io_deq_bits_id;
  wire  _T_968_valid;
  wire  _T_968_bits_id;
  reg [2:0] _T_989_0;
  reg [31:0] _RAND_9;
  reg [2:0] _T_989_1;
  reg [31:0] _RAND_10;
  wire [2:0] _GEN_12;
  wire [2:0] _GEN_13;
  wire  _T_1006;
  wire [1:0] _T_1009;
  wire  _T_1011;
  wire  _T_1012;
  wire  _T_1013;
  wire  _T_1014;
  wire [3:0] _T_1016;
  wire [2:0] _T_1017;
  wire [2:0] _GEN_14;
  wire  _T_1019;
  wire [3:0] _T_1021;
  wire [2:0] _T_1022;
  wire [2:0] _GEN_15;
  wire  _T_1023;
  wire  _T_1024;
  Queue_39 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_last(Queue_io_enq_bits_last),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_last(Queue_io_deq_bits_last)
  );
  Queue_40 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id)
  );
  assign io_in_0_aw_ready = _T_615;
  assign io_in_0_w_ready = _T_616;
  assign io_in_0_b_valid = _T_1023;
  assign io_in_0_b_bits_id = _T_968_bits_id;
  assign io_in_0_ar_ready = _T_866;
  assign io_in_0_r_valid = _T_958_valid;
  assign io_in_0_r_bits_id = _T_958_bits_id;
  assign io_in_0_r_bits_last = _T_958_bits_last;
  assign io_out_0_a_valid = _T_877;
  assign io_out_0_a_bits_opcode = _T_906;
  assign io_out_0_a_bits_param = _T_905;
  assign io_out_0_a_bits_size = _T_904;
  assign io_out_0_a_bits_source = _T_903;
  assign io_out_0_a_bits_address = _T_902;
  assign io_out_0_a_bits_mask = _T_901;
  assign io_out_0_a_bits_data = _T_900;
  assign io_out_0_d_ready = _T_947;
  assign _T_95 = {io_in_0_ar_bits_len,8'hff};
  assign _GEN_16 = {{7'd0}, _T_95};
  assign _T_96 = _GEN_16 << io_in_0_ar_bits_size;
  assign _T_97 = _T_96[22:8];
  assign _GEN_17 = {{1'd0}, _T_97};
  assign _T_98 = _GEN_17 << 1;
  assign _T_100 = _T_98 | 16'h1;
  assign _T_102 = {1'h0,_T_97};
  assign _T_103 = ~ _T_102;
  assign _T_104 = _T_100 & _T_103;
  assign _T_105 = _T_104[15:8];
  assign _T_106 = _T_104[7:0];
  assign _T_108 = _T_105 != 8'h0;
  assign _T_109 = _T_105 | _T_106;
  assign _T_110 = _T_109[7:4];
  assign _T_111 = _T_109[3:0];
  assign _T_113 = _T_110 != 4'h0;
  assign _T_114 = _T_110 | _T_111;
  assign _T_115 = _T_114[3:2];
  assign _T_116 = _T_114[1:0];
  assign _T_118 = _T_115 != 2'h0;
  assign _T_119 = _T_115 | _T_116;
  assign _T_120 = _T_119[1];
  assign _T_121 = {_T_118,_T_120};
  assign _T_122 = {_T_113,_T_121};
  assign _T_123 = {_T_108,_T_122};
  assign _T_128 = _T_123 <= 4'hc;
  assign _T_132 = io_in_0_ar_bits_addr ^ 32'h3000;
  assign _T_133 = {1'b0,$signed(_T_132)};
  assign _T_135 = $signed(_T_133) & $signed(-33'sh1000);
  assign _T_136 = $signed(_T_135);
  assign _T_138 = $signed(_T_136) == $signed(33'sh0);
  assign _T_139 = _T_128 & _T_138;
  assign _T_144 = _T_123 <= 4'h6;
  assign _T_148 = io_in_0_ar_bits_addr ^ 32'hc000000;
  assign _T_149 = {1'b0,$signed(_T_148)};
  assign _T_151 = $signed(_T_149) & $signed(-33'sh4000000);
  assign _T_152 = $signed(_T_151);
  assign _T_154 = $signed(_T_152) == $signed(33'sh0);
  assign _T_156 = io_in_0_ar_bits_addr ^ 32'h2000000;
  assign _T_157 = {1'b0,$signed(_T_156)};
  assign _T_159 = $signed(_T_157) & $signed(-33'sh10000);
  assign _T_160 = $signed(_T_159);
  assign _T_162 = $signed(_T_160) == $signed(33'sh0);
  assign _T_165 = {1'b0,$signed(io_in_0_ar_bits_addr)};
  assign _T_167 = $signed(_T_165) & $signed(-33'sh1000);
  assign _T_168 = $signed(_T_167);
  assign _T_170 = $signed(_T_168) == $signed(33'sh0);
  assign _T_172 = io_in_0_ar_bits_addr ^ 32'h10000;
  assign _T_173 = {1'b0,$signed(_T_172)};
  assign _T_175 = $signed(_T_173) & $signed(-33'sh10000);
  assign _T_176 = $signed(_T_175);
  assign _T_178 = $signed(_T_176) == $signed(33'sh0);
  assign _T_180 = io_in_0_ar_bits_addr ^ 32'h80000000;
  assign _T_181 = {1'b0,$signed(_T_180)};
  assign _T_183 = $signed(_T_181) & $signed(-33'sh4000);
  assign _T_184 = $signed(_T_183);
  assign _T_186 = $signed(_T_184) == $signed(33'sh0);
  assign _T_188 = io_in_0_ar_bits_addr ^ 32'h60000000;
  assign _T_189 = {1'b0,$signed(_T_188)};
  assign _T_191 = $signed(_T_189) & $signed(-33'sh20000000);
  assign _T_192 = $signed(_T_191);
  assign _T_194 = $signed(_T_192) == $signed(33'sh0);
  assign _T_195 = _T_154 | _T_162;
  assign _T_196 = _T_195 | _T_170;
  assign _T_197 = _T_196 | _T_178;
  assign _T_198 = _T_197 | _T_186;
  assign _T_199 = _T_198 | _T_194;
  assign _T_200 = _T_144 & _T_199;
  assign _T_203 = _T_139 | _T_200;
  assign _T_205 = io_in_0_ar_bits_addr[2:0];
  assign _GEN_18 = {{11'd0}, _T_205};
  assign _T_206 = 14'h3000 | _GEN_18;
  assign _T_207 = _T_203 ? io_in_0_ar_bits_addr : {{18'd0}, _T_206};
  assign _GEN_4 = io_in_0_ar_bits_id ? _T_225_1 : _T_225_0;
  assign _T_239 = _GEN_4[1:0];
  assign _T_241 = {io_in_0_ar_bits_id,_T_239};
  assign _T_242 = {_T_241,1'h0};
  assign _T_244 = io_in_0_ar_valid == 1'h0;
  assign _T_247 = 30'h7fff << _T_123;
  assign _T_248 = _T_247[14:0];
  assign _T_249 = ~ _T_248;
  assign _T_250 = _T_97 == _T_249;
  assign _T_251 = _T_244 | _T_250;
  assign _T_252 = _T_251 | reset;
  assign _T_254 = _T_252 == 1'h0;
  assign _T_339 = _T_123[1:0];
  assign _T_341 = 4'h1 << _T_339;
  assign _T_342 = _T_341[2:0];
  assign _T_344 = _T_342 | 3'h1;
  assign _T_346 = _T_123 >= 4'h3;
  assign _T_348 = _T_344[2];
  assign _T_349 = _T_207[2];
  assign _T_351 = _T_349 == 1'h0;
  assign _T_353 = _T_348 & _T_351;
  assign _T_354 = _T_346 | _T_353;
  assign _T_356 = _T_348 & _T_349;
  assign _T_357 = _T_346 | _T_356;
  assign _T_358 = _T_344[1];
  assign _T_359 = _T_207[1];
  assign _T_361 = _T_359 == 1'h0;
  assign _T_362 = _T_351 & _T_361;
  assign _T_363 = _T_358 & _T_362;
  assign _T_364 = _T_354 | _T_363;
  assign _T_365 = _T_351 & _T_359;
  assign _T_366 = _T_358 & _T_365;
  assign _T_367 = _T_354 | _T_366;
  assign _T_368 = _T_349 & _T_361;
  assign _T_369 = _T_358 & _T_368;
  assign _T_370 = _T_357 | _T_369;
  assign _T_371 = _T_349 & _T_359;
  assign _T_372 = _T_358 & _T_371;
  assign _T_373 = _T_357 | _T_372;
  assign _T_374 = _T_344[0];
  assign _T_375 = _T_207[0];
  assign _T_377 = _T_375 == 1'h0;
  assign _T_378 = _T_362 & _T_377;
  assign _T_379 = _T_374 & _T_378;
  assign _T_380 = _T_364 | _T_379;
  assign _T_381 = _T_362 & _T_375;
  assign _T_382 = _T_374 & _T_381;
  assign _T_383 = _T_364 | _T_382;
  assign _T_384 = _T_365 & _T_377;
  assign _T_385 = _T_374 & _T_384;
  assign _T_386 = _T_367 | _T_385;
  assign _T_387 = _T_365 & _T_375;
  assign _T_388 = _T_374 & _T_387;
  assign _T_389 = _T_367 | _T_388;
  assign _T_390 = _T_368 & _T_377;
  assign _T_391 = _T_374 & _T_390;
  assign _T_392 = _T_370 | _T_391;
  assign _T_393 = _T_368 & _T_375;
  assign _T_394 = _T_374 & _T_393;
  assign _T_395 = _T_370 | _T_394;
  assign _T_396 = _T_371 & _T_377;
  assign _T_397 = _T_374 & _T_396;
  assign _T_398 = _T_373 | _T_397;
  assign _T_399 = _T_371 & _T_375;
  assign _T_400 = _T_374 & _T_399;
  assign _T_401 = _T_373 | _T_400;
  assign _T_402 = {_T_383,_T_380};
  assign _T_403 = {_T_389,_T_386};
  assign _T_404 = {_T_403,_T_402};
  assign _T_405 = {_T_395,_T_392};
  assign _T_406 = {_T_401,_T_398};
  assign _T_407 = {_T_406,_T_405};
  assign _T_408 = {_T_407,_T_404};
  assign _T_412 = 2'h1 << io_in_0_ar_bits_id;
  assign _T_414 = _T_412[0];
  assign _T_415 = _T_412[1];
  assign _T_416 = io_in_0_ar_ready & io_in_0_ar_valid;
  assign _T_417 = _T_416 & _T_414;
  assign _T_419 = _T_225_0 + 3'h1;
  assign _T_420 = _T_419[2:0];
  assign _GEN_5 = _T_417 ? _T_420 : _T_225_0;
  assign _T_422 = _T_416 & _T_415;
  assign _T_424 = _T_225_1 + 3'h1;
  assign _T_425 = _T_424[2:0];
  assign _GEN_6 = _T_422 ? _T_425 : _T_225_1;
  assign _T_431 = {io_in_0_aw_bits_len,8'hff};
  assign _GEN_19 = {{7'd0}, _T_431};
  assign _T_432 = _GEN_19 << io_in_0_aw_bits_size;
  assign _T_433 = _T_432[22:8];
  assign _GEN_20 = {{1'd0}, _T_433};
  assign _T_434 = _GEN_20 << 1;
  assign _T_436 = _T_434 | 16'h1;
  assign _T_438 = {1'h0,_T_433};
  assign _T_439 = ~ _T_438;
  assign _T_440 = _T_436 & _T_439;
  assign _T_441 = _T_440[15:8];
  assign _T_442 = _T_440[7:0];
  assign _T_444 = _T_441 != 8'h0;
  assign _T_445 = _T_441 | _T_442;
  assign _T_446 = _T_445[7:4];
  assign _T_447 = _T_445[3:0];
  assign _T_449 = _T_446 != 4'h0;
  assign _T_450 = _T_446 | _T_447;
  assign _T_451 = _T_450[3:2];
  assign _T_452 = _T_450[1:0];
  assign _T_454 = _T_451 != 2'h0;
  assign _T_455 = _T_451 | _T_452;
  assign _T_456 = _T_455[1];
  assign _T_457 = {_T_454,_T_456};
  assign _T_458 = {_T_449,_T_457};
  assign _T_459 = {_T_444,_T_458};
  assign _T_464 = _T_459 <= 4'hc;
  assign _T_468 = io_in_0_aw_bits_addr ^ 32'h3000;
  assign _T_469 = {1'b0,$signed(_T_468)};
  assign _T_471 = $signed(_T_469) & $signed(-33'sh1000);
  assign _T_472 = $signed(_T_471);
  assign _T_474 = $signed(_T_472) == $signed(33'sh0);
  assign _T_475 = _T_464 & _T_474;
  assign _T_480 = _T_459 <= 4'h6;
  assign _T_484 = io_in_0_aw_bits_addr ^ 32'hc000000;
  assign _T_485 = {1'b0,$signed(_T_484)};
  assign _T_487 = $signed(_T_485) & $signed(-33'sh4000000);
  assign _T_488 = $signed(_T_487);
  assign _T_490 = $signed(_T_488) == $signed(33'sh0);
  assign _T_492 = io_in_0_aw_bits_addr ^ 32'h2000000;
  assign _T_493 = {1'b0,$signed(_T_492)};
  assign _T_495 = $signed(_T_493) & $signed(-33'sh10000);
  assign _T_496 = $signed(_T_495);
  assign _T_498 = $signed(_T_496) == $signed(33'sh0);
  assign _T_501 = {1'b0,$signed(io_in_0_aw_bits_addr)};
  assign _T_503 = $signed(_T_501) & $signed(-33'sh1000);
  assign _T_504 = $signed(_T_503);
  assign _T_506 = $signed(_T_504) == $signed(33'sh0);
  assign _T_508 = io_in_0_aw_bits_addr ^ 32'h80000000;
  assign _T_509 = {1'b0,$signed(_T_508)};
  assign _T_511 = $signed(_T_509) & $signed(-33'sh4000);
  assign _T_512 = $signed(_T_511);
  assign _T_514 = $signed(_T_512) == $signed(33'sh0);
  assign _T_515 = _T_490 | _T_498;
  assign _T_516 = _T_515 | _T_506;
  assign _T_517 = _T_516 | _T_514;
  assign _T_518 = _T_480 & _T_517;
  assign _T_523 = _T_459 <= 4'h8;
  assign _T_527 = io_in_0_aw_bits_addr ^ 32'h60000000;
  assign _T_528 = {1'b0,$signed(_T_527)};
  assign _T_530 = $signed(_T_528) & $signed(-33'sh20000000);
  assign _T_531 = $signed(_T_530);
  assign _T_533 = $signed(_T_531) == $signed(33'sh0);
  assign _T_534 = _T_523 & _T_533;
  assign _T_549 = _T_475 | _T_518;
  assign _T_550 = _T_549 | _T_534;
  assign _T_553 = io_in_0_aw_bits_addr[2:0];
  assign _GEN_21 = {{11'd0}, _T_553};
  assign _T_554 = 14'h3000 | _GEN_21;
  assign _T_555 = _T_550 ? io_in_0_aw_bits_addr : {{18'd0}, _T_554};
  assign _GEN_7 = io_in_0_aw_bits_id ? _T_573_1 : _T_573_0;
  assign _T_587 = _GEN_7[1:0];
  assign _T_589 = {io_in_0_aw_bits_id,_T_587};
  assign _T_590 = {_T_589,1'h1};
  assign _T_592 = io_in_0_aw_valid == 1'h0;
  assign _T_595 = 30'h7fff << _T_459;
  assign _T_596 = _T_595[14:0];
  assign _T_597 = ~ _T_596;
  assign _T_598 = _T_433 == _T_597;
  assign _T_599 = _T_592 | _T_598;
  assign _T_600 = _T_599 | reset;
  assign _T_602 = _T_600 == 1'h0;
  assign _T_606 = io_in_0_aw_bits_len == 8'h0;
  assign _T_607 = _T_592 | _T_606;
  assign _T_609 = io_in_0_aw_bits_size == 3'h3;
  assign _T_610 = _T_607 | _T_609;
  assign _T_611 = _T_610 | reset;
  assign _T_613 = _T_611 == 1'h0;
  assign _T_614 = _T_867 & io_in_0_w_valid;
  assign _T_615 = _T_614 & io_in_0_w_bits_last;
  assign _T_616 = _T_867 & io_in_0_aw_valid;
  assign _T_617 = io_in_0_aw_valid & io_in_0_w_valid;
  assign _T_716 = 2'h1 << io_in_0_aw_bits_id;
  assign _T_718 = _T_716[0];
  assign _T_719 = _T_716[1];
  assign _T_720 = io_in_0_aw_ready & io_in_0_aw_valid;
  assign _T_721 = _T_720 & _T_718;
  assign _T_723 = _T_573_0 + 3'h1;
  assign _T_724 = _T_723[2:0];
  assign _GEN_8 = _T_721 ? _T_724 : _T_573_0;
  assign _T_726 = _T_720 & _T_719;
  assign _T_728 = _T_573_1 + 3'h1;
  assign _T_729 = _T_728[2:0];
  assign _GEN_9 = _T_726 ? _T_729 : _T_573_1;
  assign _T_735 = _T_733 == 8'h0;
  assign _T_736 = _T_735 & io_out_0_a_ready;
  assign _T_737 = {_T_617,io_in_0_ar_valid};
  assign _T_739 = _T_737 == _T_737;
  assign _T_740 = _T_739 | reset;
  assign _T_742 = _T_740 == 1'h0;
  assign _T_747 = ~ _T_746;
  assign _T_748 = _T_737 & _T_747;
  assign _T_749 = {_T_748,_T_737};
  assign _T_750 = _T_749[3:1];
  assign _GEN_22 = {{1'd0}, _T_750};
  assign _T_751 = _T_749 | _GEN_22;
  assign _T_753 = _T_751[3:1];
  assign _GEN_23 = {{2'd0}, _T_746};
  assign _T_754 = _GEN_23 << 2;
  assign _GEN_24 = {{1'd0}, _T_753};
  assign _T_755 = _GEN_24 | _T_754;
  assign _T_756 = _T_755[3:2];
  assign _T_757 = _T_755[1:0];
  assign _T_758 = _T_756 & _T_757;
  assign _T_759 = ~ _T_758;
  assign _T_761 = _T_737 != 2'h0;
  assign _T_762 = _T_736 & _T_761;
  assign _T_763 = _T_759 & _T_737;
  assign _GEN_25 = {{1'd0}, _T_763};
  assign _T_764 = _GEN_25 << 1;
  assign _T_765 = _T_764[1:0];
  assign _T_766 = _T_763 | _T_765;
  assign _GEN_10 = _T_762 ? _T_766 : _T_746;
  assign _T_769 = _T_759[0];
  assign _T_770 = _T_759[1];
  assign _T_778 = _T_769 & io_in_0_ar_valid;
  assign _T_779 = _T_770 & _T_617;
  assign _T_789 = _T_778 | _T_779;
  assign _T_793 = _T_778 == 1'h0;
  assign _T_798 = _T_779 == 1'h0;
  assign _T_799 = _T_793 | _T_798;
  assign _T_801 = _T_799 | reset;
  assign _T_803 = _T_801 == 1'h0;
  assign _T_804 = io_in_0_ar_valid | _T_617;
  assign _T_806 = _T_804 == 1'h0;
  assign _T_808 = _T_806 | _T_789;
  assign _T_809 = _T_808 | reset;
  assign _T_811 = _T_809 == 1'h0;
  assign _T_815 = _T_779 ? io_in_0_aw_bits_len : 8'h0;
  assign _T_817 = io_out_0_a_ready & io_out_0_a_valid;
  assign _GEN_26 = {{7'd0}, _T_817};
  assign _T_818 = _T_733 - _GEN_26;
  assign _T_819 = $unsigned(_T_818);
  assign _T_820 = _T_819[7:0];
  assign _T_821 = _T_736 ? _T_815 : _T_820;
  assign _T_850_0 = _T_735 ? _T_778 : _T_839_0;
  assign _T_850_1 = _T_735 ? _T_779 : _T_839_1;
  assign _T_858_0 = _T_735 ? _T_769 : _T_839_0;
  assign _T_858_1 = _T_735 ? _T_770 : _T_839_1;
  assign _T_866 = io_out_0_a_ready & _T_858_0;
  assign _T_867 = io_out_0_a_ready & _T_858_1;
  assign _T_871 = _T_839_0 ? io_in_0_ar_valid : 1'h0;
  assign _T_873 = _T_839_1 ? _T_617 : 1'h0;
  assign _T_874 = _T_871 | _T_873;
  assign _T_877 = _T_735 ? _T_804 : _T_874;
  assign _T_879 = {_T_207,_T_408};
  assign _T_880 = {_T_879,64'h0};
  assign _T_881 = {_T_123,_T_242};
  assign _T_883 = {6'h20,_T_881};
  assign _T_884 = {_T_883,_T_880};
  assign _T_886 = _T_850_0 ? _T_884 : 118'h0;
  assign _T_887 = {_T_555,io_in_0_w_bits_strb};
  assign _T_888 = {_T_887,io_in_0_w_bits_data};
  assign _T_889 = {_T_459,_T_590};
  assign _T_891 = {6'h8,_T_889};
  assign _T_892 = {_T_891,_T_888};
  assign _T_894 = _T_850_1 ? _T_892 : 118'h0;
  assign _T_895 = _T_886 | _T_894;
  assign _T_900 = _T_895[63:0];
  assign _T_901 = _T_895[71:64];
  assign _T_902 = _T_895[103:72];
  assign _T_903 = _T_895[107:104];
  assign _T_904 = _T_895[111:108];
  assign _T_905 = _T_895[114:112];
  assign _T_906 = _T_895[117:115];
  assign _T_907_ready = Queue_1_io_enq_ready;
  assign _T_911_ready = Queue_io_enq_ready;
  assign _T_918 = io_out_0_d_bits_opcode[0];
  assign _T_919 = io_out_0_d_ready & io_out_0_d_valid;
  assign _T_922 = 27'hfff << io_out_0_d_bits_size;
  assign _T_923 = _T_922[11:0];
  assign _T_924 = ~ _T_923;
  assign _T_925 = _T_924[11:3];
  assign _T_928 = _T_918 ? _T_925 : 9'h0;
  assign _T_933 = _T_931 - 9'h1;
  assign _T_934 = $unsigned(_T_933);
  assign _T_935 = _T_934[8:0];
  assign _T_937 = _T_931 == 9'h0;
  assign _T_939 = _T_931 == 9'h1;
  assign _T_941 = _T_928 == 9'h0;
  assign _T_942 = _T_939 | _T_941;
  assign _T_946 = _T_937 ? _T_928 : _T_935;
  assign _GEN_11 = _T_919 ? _T_946 : _T_931;
  assign _T_947 = _T_918 ? _T_911_ready : _T_907_ready;
  assign _T_948 = io_out_0_d_valid & _T_918;
  assign _T_950 = _T_918 == 1'h0;
  assign _T_951 = io_out_0_d_valid & _T_950;
  assign _T_952 = io_out_0_d_bits_source[3:3];
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = _T_948;
  assign Queue_io_enq_bits_id = _T_952;
  assign Queue_io_enq_bits_last = _T_942;
  assign Queue_io_deq_ready = io_in_0_r_ready;
  assign _T_958_valid = Queue_io_deq_valid;
  assign _T_958_bits_id = Queue_io_deq_bits_id;
  assign _T_958_bits_last = Queue_io_deq_bits_last;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = _T_951;
  assign Queue_1_io_enq_bits_id = _T_952;
  assign Queue_1_io_deq_ready = _T_1024;
  assign _T_968_valid = Queue_1_io_deq_valid;
  assign _T_968_bits_id = Queue_1_io_deq_bits_id;
  assign _GEN_12 = io_in_0_b_bits_id ? _T_989_1 : _T_989_0;
  assign _GEN_13 = io_in_0_b_bits_id ? _T_573_1 : _T_573_0;
  assign _T_1006 = _GEN_12 != _GEN_13;
  assign _T_1009 = 2'h1 << io_in_0_b_bits_id;
  assign _T_1011 = _T_1009[0];
  assign _T_1012 = _T_1009[1];
  assign _T_1013 = io_in_0_b_ready & io_in_0_b_valid;
  assign _T_1014 = _T_1013 & _T_1011;
  assign _T_1016 = _T_989_0 + 3'h1;
  assign _T_1017 = _T_1016[2:0];
  assign _GEN_14 = _T_1014 ? _T_1017 : _T_989_0;
  assign _T_1019 = _T_1013 & _T_1012;
  assign _T_1021 = _T_989_1 + 3'h1;
  assign _T_1022 = _T_1021[2:0];
  assign _GEN_15 = _T_1019 ? _T_1022 : _T_989_1;
  assign _T_1023 = _T_968_valid & _T_1006;
  assign _T_1024 = io_in_0_b_ready & _T_1006;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_225_0 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_225_1 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_573_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_573_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_733 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_746 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_839_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_839_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_931 = _RAND_8[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_989_0 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_989_1 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225_0 <= 3'h0;
    end else begin
      if (_T_417) begin
        _T_225_0 <= _T_420;
      end
    end
    if (reset) begin
      _T_225_1 <= 3'h0;
    end else begin
      if (_T_422) begin
        _T_225_1 <= _T_425;
      end
    end
    if (reset) begin
      _T_573_0 <= 3'h0;
    end else begin
      if (_T_721) begin
        _T_573_0 <= _T_724;
      end
    end
    if (reset) begin
      _T_573_1 <= 3'h0;
    end else begin
      if (_T_726) begin
        _T_573_1 <= _T_729;
      end
    end
    if (reset) begin
      _T_733 <= 8'h0;
    end else begin
      if (_T_736) begin
        if (_T_779) begin
          _T_733 <= io_in_0_aw_bits_len;
        end else begin
          _T_733 <= 8'h0;
        end
      end else begin
        _T_733 <= _T_820;
      end
    end
    if (reset) begin
      _T_746 <= 2'h3;
    end else begin
      if (_T_762) begin
        _T_746 <= _T_766;
      end
    end
    if (reset) begin
      _T_839_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        _T_839_0 <= _T_778;
      end
    end
    if (reset) begin
      _T_839_1 <= 1'h0;
    end else begin
      if (_T_735) begin
        _T_839_1 <= _T_779;
      end
    end
    if (reset) begin
      _T_931 <= 9'h0;
    end else begin
      if (_T_919) begin
        if (_T_937) begin
          if (_T_918) begin
            _T_931 <= _T_925;
          end else begin
            _T_931 <= 9'h0;
          end
        end else begin
          _T_931 <= _T_935;
        end
      end
    end
    if (reset) begin
      _T_989_0 <= 3'h0;
    end else begin
      if (_T_1014) begin
        _T_989_0 <= _T_1017;
      end
    end
    if (reset) begin
      _T_989_1 <= 3'h0;
    end else begin
      if (_T_1019) begin
        _T_989_1 <= _T_1022;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_254) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:82 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_254) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_602) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:100 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_602) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_613) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToTL.scala:101 assert (!in.aw.valid || in.aw.bits.len === UInt(0) || in.aw.bits.size === UInt(log2Ceil(beatBytes))) // because aligned\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_613) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_742) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:19 assert (valid === valids)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_742) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_803) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_803) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_811) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_811) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Repeater_6(
  input         clock,
  input         reset,
  input         io_repeat,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [2:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [3:0]  io_enq_bits_source,
  input  [31:0] io_enq_bits_address,
  input  [7:0]  io_enq_bits_mask,
  input  [63:0] io_enq_bits_data,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [2:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [3:0]  io_deq_bits_source,
  output [31:0] io_deq_bits_address,
  output [7:0]  io_deq_bits_mask,
  output [63:0] io_deq_bits_data
);
  reg  full;
  reg [31:0] _RAND_0;
  reg [2:0] saved_opcode;
  reg [31:0] _RAND_1;
  reg [2:0] saved_param;
  reg [31:0] _RAND_2;
  reg [3:0] saved_size;
  reg [31:0] _RAND_3;
  reg [3:0] saved_source;
  reg [31:0] _RAND_4;
  reg [31:0] saved_address;
  reg [31:0] _RAND_5;
  reg [7:0] saved_mask;
  reg [31:0] _RAND_6;
  reg [63:0] saved_data;
  reg [63:0] _RAND_7;
  wire  _T_16;
  wire  _T_18;
  wire  _T_19;
  wire [2:0] _T_20_opcode;
  wire [2:0] _T_20_param;
  wire [3:0] _T_20_size;
  wire [3:0] _T_20_source;
  wire [31:0] _T_20_address;
  wire [7:0] _T_20_mask;
  wire [63:0] _T_20_data;
  wire  _T_21;
  wire  _T_22;
  wire  _GEN_0;
  wire [2:0] _GEN_1;
  wire [2:0] _GEN_2;
  wire [3:0] _GEN_3;
  wire [3:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [7:0] _GEN_6;
  wire [63:0] _GEN_7;
  wire  _T_24;
  wire  _T_26;
  wire  _T_27;
  wire  _GEN_8;
  assign io_enq_ready = _T_19;
  assign io_deq_valid = _T_16;
  assign io_deq_bits_opcode = _T_20_opcode;
  assign io_deq_bits_param = _T_20_param;
  assign io_deq_bits_size = _T_20_size;
  assign io_deq_bits_source = _T_20_source;
  assign io_deq_bits_address = _T_20_address;
  assign io_deq_bits_mask = _T_20_mask;
  assign io_deq_bits_data = _T_20_data;
  assign _T_16 = io_enq_valid | full;
  assign _T_18 = full == 1'h0;
  assign _T_19 = io_deq_ready & _T_18;
  assign _T_20_opcode = full ? saved_opcode : io_enq_bits_opcode;
  assign _T_20_param = full ? saved_param : io_enq_bits_param;
  assign _T_20_size = full ? saved_size : io_enq_bits_size;
  assign _T_20_source = full ? saved_source : io_enq_bits_source;
  assign _T_20_address = full ? saved_address : io_enq_bits_address;
  assign _T_20_mask = full ? saved_mask : io_enq_bits_mask;
  assign _T_20_data = full ? saved_data : io_enq_bits_data;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_22 = _T_21 & io_repeat;
  assign _GEN_0 = _T_22 ? 1'h1 : full;
  assign _GEN_1 = _T_22 ? io_enq_bits_opcode : saved_opcode;
  assign _GEN_2 = _T_22 ? io_enq_bits_param : saved_param;
  assign _GEN_3 = _T_22 ? io_enq_bits_size : saved_size;
  assign _GEN_4 = _T_22 ? io_enq_bits_source : saved_source;
  assign _GEN_5 = _T_22 ? io_enq_bits_address : saved_address;
  assign _GEN_6 = _T_22 ? io_enq_bits_mask : saved_mask;
  assign _GEN_7 = _T_22 ? io_enq_bits_data : saved_data;
  assign _T_24 = io_deq_ready & io_deq_valid;
  assign _T_26 = io_repeat == 1'h0;
  assign _T_27 = _T_24 & _T_26;
  assign _GEN_8 = _T_27 ? 1'h0 : _GEN_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  saved_opcode = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  saved_param = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  saved_size = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  saved_source = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  saved_address = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  saved_mask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{$random}};
  saved_data = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      full <= 1'h0;
    end else begin
      if (_T_27) begin
        full <= 1'h0;
      end else begin
        if (_T_22) begin
          full <= 1'h1;
        end
      end
    end
    if (_T_22) begin
      saved_opcode <= io_enq_bits_opcode;
    end
    if (_T_22) begin
      saved_param <= io_enq_bits_param;
    end
    if (_T_22) begin
      saved_size <= io_enq_bits_size;
    end
    if (_T_22) begin
      saved_source <= io_enq_bits_source;
    end
    if (_T_22) begin
      saved_address <= io_enq_bits_address;
    end
    if (_T_22) begin
      saved_mask <= io_enq_bits_mask;
    end
    if (_T_22) begin
      saved_data <= io_enq_bits_data;
    end
  end
endmodule
module TLWidthWidget_2(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [2:0]  io_in_0_a_bits_param,
  input  [3:0]  io_in_0_a_bits_size,
  input  [3:0]  io_in_0_a_bits_source,
  input  [31:0] io_in_0_a_bits_address,
  input  [7:0]  io_in_0_a_bits_mask,
  input  [63:0] io_in_0_a_bits_data,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [3:0]  io_in_0_d_bits_size,
  output [3:0]  io_in_0_d_bits_source,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [2:0]  io_out_0_a_bits_param,
  output [3:0]  io_out_0_a_bits_size,
  output [3:0]  io_out_0_a_bits_source,
  output [31:0] io_out_0_a_bits_address,
  output [3:0]  io_out_0_a_bits_mask,
  output [31:0] io_out_0_a_bits_data,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [3:0]  io_out_0_d_bits_size,
  input  [3:0]  io_out_0_d_bits_source
);
  wire  Repeater_clock;
  wire  Repeater_reset;
  wire  Repeater_io_repeat;
  wire  Repeater_io_enq_ready;
  wire  Repeater_io_enq_valid;
  wire [2:0] Repeater_io_enq_bits_opcode;
  wire [2:0] Repeater_io_enq_bits_param;
  wire [3:0] Repeater_io_enq_bits_size;
  wire [3:0] Repeater_io_enq_bits_source;
  wire [31:0] Repeater_io_enq_bits_address;
  wire [7:0] Repeater_io_enq_bits_mask;
  wire [63:0] Repeater_io_enq_bits_data;
  wire  Repeater_io_deq_ready;
  wire  Repeater_io_deq_valid;
  wire [2:0] Repeater_io_deq_bits_opcode;
  wire [2:0] Repeater_io_deq_bits_param;
  wire [3:0] Repeater_io_deq_bits_size;
  wire [3:0] Repeater_io_deq_bits_source;
  wire [31:0] Repeater_io_deq_bits_address;
  wire [7:0] Repeater_io_deq_bits_mask;
  wire [63:0] Repeater_io_deq_bits_data;
  wire  _T_92_valid;
  wire [2:0] _T_92_bits_opcode;
  wire [2:0] _T_92_bits_param;
  wire [3:0] _T_92_bits_size;
  wire [3:0] _T_92_bits_source;
  wire [31:0] _T_92_bits_address;
  wire [7:0] _T_92_bits_mask;
  wire [31:0] _T_96;
  wire [31:0] _T_97;
  wire [63:0] _T_98;
  wire  _T_99;
  wire  _T_101;
  wire [17:0] _T_104;
  wire [2:0] _T_105;
  wire [2:0] _T_106;
  wire  _T_107;
  reg  _T_110;
  reg [31:0] _RAND_0;
  wire  _T_113;
  wire  _T_115;
  wire  _T_116;
  wire  _T_117;
  wire [1:0] _T_119;
  wire  _T_120;
  wire  _GEN_2;
  wire  _GEN_3;
  wire  _T_122;
  wire  _T_123;
  wire [31:0] _T_124;
  wire [31:0] _T_125;
  wire [31:0] _GEN_4;
  wire [3:0] _T_134;
  wire [3:0] _T_135;
  wire [3:0] _GEN_5;
  wire  _T_145;
  wire  _T_146;
  wire [17:0] _T_149;
  wire [2:0] _T_150;
  wire [2:0] _T_151;
  wire  _T_152;
  reg  _T_155;
  reg [31:0] _RAND_1;
  wire  _T_158;
  wire  _T_160;
  wire  _T_161;
  wire  _T_176;
  wire [1:0] _T_178;
  wire  _T_179;
  wire  _GEN_6;
  wire  _GEN_7;
  wire  _T_182;
  wire  _T_183;
  wire  _T_184;
  Repeater_6 Repeater (
    .clock(Repeater_clock),
    .reset(Repeater_reset),
    .io_repeat(Repeater_io_repeat),
    .io_enq_ready(Repeater_io_enq_ready),
    .io_enq_valid(Repeater_io_enq_valid),
    .io_enq_bits_opcode(Repeater_io_enq_bits_opcode),
    .io_enq_bits_param(Repeater_io_enq_bits_param),
    .io_enq_bits_size(Repeater_io_enq_bits_size),
    .io_enq_bits_source(Repeater_io_enq_bits_source),
    .io_enq_bits_address(Repeater_io_enq_bits_address),
    .io_enq_bits_mask(Repeater_io_enq_bits_mask),
    .io_enq_bits_data(Repeater_io_enq_bits_data),
    .io_deq_ready(Repeater_io_deq_ready),
    .io_deq_valid(Repeater_io_deq_valid),
    .io_deq_bits_opcode(Repeater_io_deq_bits_opcode),
    .io_deq_bits_param(Repeater_io_deq_bits_param),
    .io_deq_bits_size(Repeater_io_deq_bits_size),
    .io_deq_bits_source(Repeater_io_deq_bits_source),
    .io_deq_bits_address(Repeater_io_deq_bits_address),
    .io_deq_bits_mask(Repeater_io_deq_bits_mask),
    .io_deq_bits_data(Repeater_io_deq_bits_data)
  );
  assign io_in_0_a_ready = Repeater_io_enq_ready;
  assign io_in_0_d_valid = _T_184;
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode;
  assign io_in_0_d_bits_size = io_out_0_d_bits_size;
  assign io_in_0_d_bits_source = io_out_0_d_bits_source;
  assign io_out_0_a_valid = _T_92_valid;
  assign io_out_0_a_bits_opcode = _T_92_bits_opcode;
  assign io_out_0_a_bits_param = _T_92_bits_param;
  assign io_out_0_a_bits_size = _T_92_bits_size;
  assign io_out_0_a_bits_source = _T_92_bits_source;
  assign io_out_0_a_bits_address = _T_92_bits_address;
  assign io_out_0_a_bits_mask = _GEN_5;
  assign io_out_0_a_bits_data = _GEN_4;
  assign io_out_0_d_ready = _T_183;
  assign Repeater_clock = clock;
  assign Repeater_reset = reset;
  assign Repeater_io_repeat = _T_145;
  assign Repeater_io_enq_valid = io_in_0_a_valid;
  assign Repeater_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Repeater_io_enq_bits_param = io_in_0_a_bits_param;
  assign Repeater_io_enq_bits_size = io_in_0_a_bits_size;
  assign Repeater_io_enq_bits_source = io_in_0_a_bits_source;
  assign Repeater_io_enq_bits_address = io_in_0_a_bits_address;
  assign Repeater_io_enq_bits_mask = io_in_0_a_bits_mask;
  assign Repeater_io_enq_bits_data = io_in_0_a_bits_data;
  assign Repeater_io_deq_ready = io_out_0_a_ready;
  assign _T_92_valid = Repeater_io_deq_valid;
  assign _T_92_bits_opcode = Repeater_io_deq_bits_opcode;
  assign _T_92_bits_param = Repeater_io_deq_bits_param;
  assign _T_92_bits_size = Repeater_io_deq_bits_size;
  assign _T_92_bits_source = Repeater_io_deq_bits_source;
  assign _T_92_bits_address = Repeater_io_deq_bits_address;
  assign _T_92_bits_mask = Repeater_io_deq_bits_mask;
  assign _T_96 = Repeater_io_deq_bits_data[63:32];
  assign _T_97 = io_in_0_a_bits_data[31:0];
  assign _T_98 = {_T_96,_T_97};
  assign _T_99 = _T_92_bits_opcode[2];
  assign _T_101 = _T_99 == 1'h0;
  assign _T_104 = 18'h7 << _T_92_bits_size;
  assign _T_105 = _T_104[2:0];
  assign _T_106 = ~ _T_105;
  assign _T_107 = _T_106[2:2];
  assign _T_113 = _T_110 == _T_107;
  assign _T_115 = _T_101 == 1'h0;
  assign _T_116 = _T_113 | _T_115;
  assign _T_117 = io_out_0_a_ready & io_out_0_a_valid;
  assign _T_119 = _T_110 + 1'h1;
  assign _T_120 = _T_119[0:0];
  assign _GEN_2 = _T_116 ? 1'h0 : _T_120;
  assign _GEN_3 = _T_117 ? _GEN_2 : _T_110;
  assign _T_122 = _T_92_bits_address[2];
  assign _T_123 = _T_122 | _T_110;
  assign _T_124 = _T_98[31:0];
  assign _T_125 = _T_98[63:32];
  assign _GEN_4 = _T_123 ? _T_125 : _T_124;
  assign _T_134 = _T_92_bits_mask[3:0];
  assign _T_135 = _T_92_bits_mask[7:4];
  assign _GEN_5 = _T_123 ? _T_135 : _T_134;
  assign _T_145 = _T_116 == 1'h0;
  assign _T_146 = io_out_0_d_bits_opcode[0];
  assign _T_149 = 18'h7 << io_out_0_d_bits_size;
  assign _T_150 = _T_149[2:0];
  assign _T_151 = ~ _T_150;
  assign _T_152 = _T_151[2:2];
  assign _T_158 = _T_155 == _T_152;
  assign _T_160 = _T_146 == 1'h0;
  assign _T_161 = _T_158 | _T_160;
  assign _T_176 = io_out_0_d_ready & io_out_0_d_valid;
  assign _T_178 = _T_155 + 1'h1;
  assign _T_179 = _T_178[0:0];
  assign _GEN_6 = _T_161 ? 1'h0 : _T_179;
  assign _GEN_7 = _T_176 ? _GEN_6 : _T_155;
  assign _T_182 = _T_161 == 1'h0;
  assign _T_183 = io_in_0_d_ready | _T_182;
  assign _T_184 = io_out_0_d_valid & _T_161;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_110 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_155 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_110 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (_T_116) begin
          _T_110 <= 1'h0;
        end else begin
          _T_110 <= _T_120;
        end
      end
    end
    if (reset) begin
      _T_155 <= 1'h0;
    end else begin
      if (_T_176) begin
        if (_T_161) begin
          _T_155 <= 1'h0;
        end else begin
          _T_155 <= _T_179;
        end
      end
    end
  end
endmodule
module TLROM_bootrom(
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [1:0]  io_in_0_a_bits_size,
  input  [9:0]  io_in_0_a_bits_source,
  input  [16:0] io_in_0_a_bits_address,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [1:0]  io_in_0_d_bits_size,
  output [9:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error
);
  wire [9:0] index;
  wire [3:0] high;
  wire  _T_2113;
  wire [31:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_7;
  wire [31:0] _GEN_8;
  wire [31:0] _GEN_9;
  wire [31:0] _GEN_10;
  wire [31:0] _GEN_11;
  wire [31:0] _GEN_12;
  wire [31:0] _GEN_13;
  wire [31:0] _GEN_14;
  wire [31:0] _GEN_15;
  wire [31:0] _GEN_16;
  wire [31:0] _GEN_17;
  wire [31:0] _GEN_18;
  wire [31:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire [31:0] _GEN_21;
  wire [31:0] _GEN_22;
  wire [31:0] _GEN_23;
  wire [31:0] _GEN_24;
  wire [31:0] _GEN_25;
  wire [31:0] _GEN_26;
  wire [31:0] _GEN_27;
  wire [31:0] _GEN_28;
  wire [31:0] _GEN_29;
  wire [31:0] _GEN_30;
  wire [31:0] _GEN_31;
  wire [31:0] _GEN_32;
  wire [31:0] _GEN_33;
  wire [31:0] _GEN_34;
  wire [31:0] _GEN_35;
  wire [31:0] _GEN_36;
  wire [31:0] _GEN_37;
  wire [31:0] _GEN_38;
  wire [31:0] _GEN_39;
  wire [31:0] _GEN_40;
  wire [31:0] _GEN_41;
  wire [31:0] _GEN_42;
  wire [31:0] _GEN_43;
  wire [31:0] _GEN_44;
  wire [31:0] _GEN_45;
  wire [31:0] _GEN_46;
  wire [31:0] _GEN_47;
  wire [31:0] _GEN_48;
  wire [31:0] _GEN_49;
  wire [31:0] _GEN_50;
  wire [31:0] _GEN_51;
  wire [31:0] _GEN_52;
  wire [31:0] _GEN_53;
  wire [31:0] _GEN_54;
  wire [31:0] _GEN_55;
  wire [31:0] _GEN_56;
  wire [31:0] _GEN_57;
  wire [31:0] _GEN_58;
  wire [31:0] _GEN_59;
  wire [31:0] _GEN_60;
  wire [31:0] _GEN_61;
  wire [31:0] _GEN_62;
  wire [31:0] _GEN_63;
  wire [31:0] _GEN_64;
  wire [31:0] _GEN_65;
  wire [31:0] _GEN_66;
  wire [31:0] _GEN_67;
  wire [31:0] _GEN_68;
  wire [31:0] _GEN_69;
  wire [31:0] _GEN_70;
  wire [31:0] _GEN_71;
  wire [31:0] _GEN_72;
  wire [31:0] _GEN_73;
  wire [31:0] _GEN_74;
  wire [31:0] _GEN_75;
  wire [31:0] _GEN_76;
  wire [31:0] _GEN_77;
  wire [31:0] _GEN_78;
  wire [31:0] _GEN_79;
  wire [31:0] _GEN_80;
  wire [31:0] _GEN_81;
  wire [31:0] _GEN_82;
  wire [31:0] _GEN_83;
  wire [31:0] _GEN_84;
  wire [31:0] _GEN_85;
  wire [31:0] _GEN_86;
  wire [31:0] _GEN_87;
  wire [31:0] _GEN_88;
  wire [31:0] _GEN_89;
  wire [31:0] _GEN_90;
  wire [31:0] _GEN_91;
  wire [31:0] _GEN_92;
  wire [31:0] _GEN_93;
  wire [31:0] _GEN_94;
  wire [31:0] _GEN_95;
  wire [31:0] _GEN_96;
  wire [31:0] _GEN_97;
  wire [31:0] _GEN_98;
  wire [31:0] _GEN_99;
  wire [31:0] _GEN_100;
  wire [31:0] _GEN_101;
  wire [31:0] _GEN_102;
  wire [31:0] _GEN_103;
  wire [31:0] _GEN_104;
  wire [31:0] _GEN_105;
  wire [31:0] _GEN_106;
  wire [31:0] _GEN_107;
  wire [31:0] _GEN_108;
  wire [31:0] _GEN_109;
  wire [31:0] _GEN_110;
  wire [31:0] _GEN_111;
  wire [31:0] _GEN_112;
  wire [31:0] _GEN_113;
  wire [31:0] _GEN_114;
  wire [31:0] _GEN_115;
  wire [31:0] _GEN_116;
  wire [31:0] _GEN_117;
  wire [31:0] _GEN_118;
  wire [31:0] _GEN_119;
  wire [31:0] _GEN_120;
  wire [31:0] _GEN_121;
  wire [31:0] _GEN_122;
  wire [31:0] _GEN_123;
  wire [31:0] _GEN_124;
  wire [31:0] _GEN_125;
  wire [31:0] _GEN_126;
  wire [31:0] _GEN_127;
  wire [31:0] _GEN_128;
  wire [31:0] _GEN_129;
  wire [31:0] _GEN_130;
  wire [31:0] _GEN_131;
  wire [31:0] _GEN_132;
  wire [31:0] _GEN_133;
  wire [31:0] _GEN_134;
  wire [31:0] _GEN_135;
  wire [31:0] _GEN_136;
  wire [31:0] _GEN_137;
  wire [31:0] _GEN_138;
  wire [31:0] _GEN_139;
  wire [31:0] _GEN_140;
  wire [31:0] _GEN_141;
  wire [31:0] _GEN_142;
  wire [31:0] _GEN_143;
  wire [31:0] _GEN_144;
  wire [31:0] _GEN_145;
  wire [31:0] _GEN_146;
  wire [31:0] _GEN_147;
  wire [31:0] _GEN_148;
  wire [31:0] _GEN_149;
  wire [31:0] _GEN_150;
  wire [31:0] _GEN_151;
  wire [31:0] _GEN_152;
  wire [31:0] _GEN_153;
  wire [31:0] _GEN_154;
  wire [31:0] _GEN_155;
  wire [31:0] _GEN_156;
  wire [31:0] _GEN_157;
  wire [31:0] _GEN_158;
  wire [31:0] _GEN_159;
  wire [31:0] _GEN_160;
  wire [31:0] _GEN_161;
  wire [31:0] _GEN_162;
  wire [31:0] _GEN_163;
  wire [31:0] _GEN_164;
  wire [31:0] _GEN_165;
  wire [31:0] _GEN_166;
  wire [31:0] _GEN_167;
  wire [31:0] _GEN_168;
  wire [31:0] _GEN_169;
  wire [31:0] _GEN_170;
  wire [31:0] _GEN_171;
  wire [31:0] _GEN_172;
  wire [31:0] _GEN_173;
  wire [31:0] _GEN_174;
  wire [31:0] _GEN_175;
  wire [31:0] _GEN_176;
  wire [31:0] _GEN_177;
  wire [31:0] _GEN_178;
  wire [31:0] _GEN_179;
  wire [31:0] _GEN_180;
  wire [31:0] _GEN_181;
  wire [31:0] _GEN_182;
  wire [31:0] _GEN_183;
  wire [31:0] _GEN_184;
  wire [31:0] _GEN_185;
  wire [31:0] _GEN_186;
  wire [31:0] _GEN_187;
  wire [31:0] _GEN_188;
  wire [31:0] _GEN_189;
  wire [31:0] _GEN_190;
  wire [31:0] _GEN_191;
  wire [31:0] _GEN_192;
  wire [31:0] _GEN_193;
  wire [31:0] _GEN_194;
  wire [31:0] _GEN_195;
  wire [31:0] _GEN_196;
  wire [31:0] _GEN_197;
  wire [31:0] _GEN_198;
  wire [31:0] _GEN_199;
  wire [31:0] _GEN_200;
  wire [31:0] _GEN_201;
  wire [31:0] _GEN_202;
  wire [31:0] _GEN_203;
  wire [31:0] _GEN_204;
  wire [31:0] _GEN_205;
  wire [31:0] _GEN_206;
  wire [31:0] _GEN_207;
  wire [31:0] _GEN_208;
  wire [31:0] _GEN_209;
  wire [31:0] _GEN_210;
  wire [31:0] _GEN_211;
  wire [31:0] _GEN_212;
  wire [31:0] _GEN_213;
  wire [31:0] _GEN_214;
  wire [31:0] _GEN_215;
  wire [31:0] _GEN_216;
  wire [31:0] _GEN_217;
  wire [31:0] _GEN_218;
  wire [31:0] _GEN_219;
  wire [31:0] _GEN_220;
  wire [31:0] _GEN_221;
  wire [31:0] _GEN_222;
  wire [31:0] _GEN_223;
  wire [31:0] _GEN_224;
  wire [31:0] _GEN_225;
  wire [31:0] _GEN_226;
  wire [31:0] _GEN_227;
  wire [31:0] _GEN_228;
  wire [31:0] _GEN_229;
  wire [31:0] _GEN_230;
  wire [31:0] _GEN_231;
  wire [31:0] _GEN_232;
  wire [31:0] _GEN_233;
  wire [31:0] _GEN_234;
  wire [31:0] _GEN_235;
  wire [31:0] _GEN_236;
  wire [31:0] _GEN_237;
  wire [31:0] _GEN_238;
  wire [31:0] _GEN_239;
  wire [31:0] _GEN_240;
  wire [31:0] _GEN_241;
  wire [31:0] _GEN_242;
  wire [31:0] _GEN_243;
  wire [31:0] _GEN_244;
  wire [31:0] _GEN_245;
  wire [31:0] _GEN_246;
  wire [31:0] _GEN_247;
  wire [31:0] _GEN_248;
  wire [31:0] _GEN_249;
  wire [31:0] _GEN_250;
  wire [31:0] _GEN_251;
  wire [31:0] _GEN_252;
  wire [31:0] _GEN_253;
  wire [31:0] _GEN_254;
  wire [31:0] _GEN_255;
  wire [31:0] _GEN_256;
  wire [31:0] _GEN_257;
  wire [31:0] _GEN_258;
  wire [31:0] _GEN_259;
  wire [31:0] _GEN_260;
  wire [31:0] _GEN_261;
  wire [31:0] _GEN_262;
  wire [31:0] _GEN_263;
  wire [31:0] _GEN_264;
  wire [31:0] _GEN_265;
  wire [31:0] _GEN_266;
  wire [31:0] _GEN_267;
  wire [31:0] _GEN_268;
  wire [31:0] _GEN_269;
  wire [31:0] _GEN_270;
  wire [31:0] _GEN_271;
  wire [31:0] _GEN_272;
  wire [31:0] _GEN_273;
  wire [31:0] _GEN_274;
  wire [31:0] _GEN_275;
  wire [31:0] _GEN_276;
  wire [31:0] _GEN_277;
  wire [31:0] _GEN_278;
  wire [31:0] _GEN_279;
  wire [31:0] _GEN_280;
  wire [31:0] _GEN_281;
  wire [31:0] _GEN_282;
  wire [31:0] _GEN_283;
  wire [31:0] _GEN_284;
  wire [31:0] _GEN_285;
  wire [31:0] _GEN_286;
  wire [31:0] _GEN_287;
  wire [31:0] _GEN_288;
  wire [31:0] _GEN_289;
  wire [31:0] _GEN_290;
  wire [31:0] _GEN_291;
  wire [31:0] _GEN_292;
  wire [31:0] _GEN_293;
  wire [31:0] _GEN_294;
  wire [31:0] _GEN_295;
  wire [31:0] _GEN_296;
  wire [31:0] _GEN_297;
  wire [31:0] _GEN_298;
  wire [31:0] _GEN_299;
  wire [31:0] _GEN_300;
  wire [31:0] _GEN_301;
  wire [31:0] _GEN_302;
  wire [31:0] _GEN_303;
  wire [31:0] _GEN_304;
  wire [31:0] _GEN_305;
  wire [31:0] _GEN_306;
  wire [31:0] _GEN_307;
  wire [31:0] _GEN_308;
  wire [31:0] _GEN_309;
  wire [31:0] _GEN_310;
  wire [31:0] _GEN_311;
  wire [31:0] _GEN_312;
  wire [31:0] _GEN_313;
  wire [31:0] _GEN_314;
  wire [31:0] _GEN_315;
  wire [31:0] _GEN_316;
  wire [31:0] _GEN_317;
  wire [31:0] _GEN_318;
  wire [31:0] _GEN_319;
  wire [31:0] _GEN_320;
  wire [31:0] _GEN_321;
  wire [31:0] _GEN_322;
  wire [31:0] _GEN_323;
  wire [31:0] _GEN_324;
  wire [31:0] _GEN_325;
  wire [31:0] _GEN_326;
  wire [31:0] _GEN_327;
  wire [31:0] _GEN_328;
  wire [31:0] _GEN_329;
  wire [31:0] _GEN_330;
  wire [31:0] _GEN_331;
  wire [31:0] _GEN_332;
  wire [31:0] _GEN_333;
  wire [31:0] _GEN_334;
  wire [31:0] _GEN_335;
  wire [31:0] _GEN_336;
  wire [31:0] _GEN_337;
  wire [31:0] _GEN_338;
  wire [31:0] _GEN_339;
  wire [31:0] _GEN_340;
  wire [31:0] _GEN_341;
  wire [31:0] _GEN_342;
  wire [31:0] _GEN_343;
  wire [31:0] _GEN_344;
  wire [31:0] _GEN_345;
  wire [31:0] _GEN_346;
  wire [31:0] _GEN_347;
  wire [31:0] _GEN_348;
  wire [31:0] _GEN_349;
  wire [31:0] _GEN_350;
  wire [31:0] _GEN_351;
  wire [31:0] _GEN_352;
  wire [31:0] _GEN_353;
  wire [31:0] _GEN_354;
  wire [31:0] _GEN_355;
  wire [31:0] _GEN_356;
  wire [31:0] _GEN_357;
  wire [31:0] _GEN_358;
  wire [31:0] _GEN_359;
  wire [31:0] _GEN_360;
  wire [31:0] _GEN_361;
  wire [31:0] _GEN_362;
  wire [31:0] _GEN_363;
  wire [31:0] _GEN_364;
  wire [31:0] _GEN_365;
  wire [31:0] _GEN_366;
  wire [31:0] _GEN_367;
  wire [31:0] _GEN_368;
  wire [31:0] _GEN_369;
  wire [31:0] _GEN_370;
  wire [31:0] _GEN_371;
  wire [31:0] _GEN_372;
  wire [31:0] _GEN_373;
  wire [31:0] _GEN_374;
  wire [31:0] _GEN_375;
  wire [31:0] _GEN_376;
  wire [31:0] _GEN_377;
  wire [31:0] _GEN_378;
  wire [31:0] _GEN_379;
  wire [31:0] _GEN_380;
  wire [31:0] _GEN_381;
  wire [31:0] _GEN_382;
  wire [31:0] _GEN_383;
  wire [31:0] _GEN_384;
  wire [31:0] _GEN_385;
  wire [31:0] _GEN_386;
  wire [31:0] _GEN_387;
  wire [31:0] _GEN_388;
  wire [31:0] _GEN_389;
  wire [31:0] _GEN_390;
  wire [31:0] _GEN_391;
  wire [31:0] _GEN_392;
  wire [31:0] _GEN_393;
  wire [31:0] _GEN_394;
  wire [31:0] _GEN_395;
  wire [31:0] _GEN_396;
  wire [31:0] _GEN_397;
  wire [31:0] _GEN_398;
  wire [31:0] _GEN_399;
  wire [31:0] _GEN_400;
  wire [31:0] _GEN_401;
  wire [31:0] _GEN_402;
  wire [31:0] _GEN_403;
  wire [31:0] _GEN_404;
  wire [31:0] _GEN_405;
  wire [31:0] _GEN_406;
  wire [31:0] _GEN_407;
  wire [31:0] _GEN_408;
  wire [31:0] _GEN_409;
  wire [31:0] _GEN_410;
  wire [31:0] _GEN_411;
  wire [31:0] _GEN_412;
  wire [31:0] _GEN_413;
  wire [31:0] _GEN_414;
  wire [31:0] _GEN_415;
  wire [31:0] _GEN_416;
  wire [31:0] _GEN_417;
  wire [31:0] _GEN_418;
  wire [31:0] _GEN_419;
  wire [31:0] _GEN_420;
  wire [31:0] _GEN_421;
  wire [31:0] _GEN_422;
  wire [31:0] _GEN_423;
  wire [31:0] _GEN_424;
  wire [31:0] _GEN_425;
  wire [31:0] _GEN_426;
  wire [31:0] _GEN_427;
  wire [31:0] _GEN_428;
  wire [31:0] _GEN_429;
  wire [31:0] _GEN_430;
  wire [31:0] _GEN_431;
  wire [31:0] _GEN_432;
  wire [31:0] _GEN_433;
  wire [31:0] _GEN_434;
  wire [31:0] _GEN_435;
  wire [31:0] _GEN_436;
  wire [31:0] _GEN_437;
  wire [31:0] _GEN_438;
  wire [31:0] _GEN_439;
  wire [31:0] _GEN_440;
  wire [31:0] _GEN_441;
  wire [31:0] _GEN_442;
  wire [31:0] _GEN_443;
  wire [31:0] _GEN_444;
  wire [31:0] _GEN_445;
  wire [31:0] _GEN_446;
  wire [31:0] _GEN_447;
  wire [31:0] _GEN_448;
  wire [31:0] _GEN_449;
  wire [31:0] _GEN_450;
  wire [31:0] _GEN_451;
  wire [31:0] _GEN_452;
  wire [31:0] _GEN_453;
  wire [31:0] _GEN_454;
  wire [31:0] _GEN_455;
  wire [31:0] _GEN_456;
  wire [31:0] _GEN_457;
  wire [31:0] _GEN_458;
  wire [31:0] _GEN_459;
  wire [31:0] _GEN_460;
  wire [31:0] _GEN_461;
  wire [31:0] _GEN_462;
  wire [31:0] _GEN_463;
  wire [31:0] _GEN_464;
  wire [31:0] _GEN_465;
  wire [31:0] _GEN_466;
  wire [31:0] _GEN_467;
  wire [31:0] _GEN_468;
  wire [31:0] _GEN_469;
  wire [31:0] _GEN_470;
  wire [31:0] _GEN_471;
  wire [31:0] _GEN_472;
  wire [31:0] _GEN_473;
  wire [31:0] _GEN_474;
  wire [31:0] _GEN_475;
  wire [31:0] _GEN_476;
  wire [31:0] _GEN_477;
  wire [31:0] _GEN_478;
  wire [31:0] _GEN_479;
  wire [31:0] _GEN_480;
  wire [31:0] _GEN_481;
  wire [31:0] _GEN_482;
  wire [31:0] _GEN_483;
  wire [31:0] _GEN_484;
  wire [31:0] _GEN_485;
  wire [31:0] _GEN_486;
  wire [31:0] _GEN_487;
  wire [31:0] _GEN_488;
  wire [31:0] _GEN_489;
  wire [31:0] _GEN_490;
  wire [31:0] _GEN_491;
  wire [31:0] _GEN_492;
  wire [31:0] _GEN_493;
  wire [31:0] _GEN_494;
  wire [31:0] _GEN_495;
  wire [31:0] _GEN_496;
  wire [31:0] _GEN_497;
  wire [31:0] _GEN_498;
  wire [31:0] _GEN_499;
  wire [31:0] _GEN_500;
  wire [31:0] _GEN_501;
  wire [31:0] _GEN_502;
  wire [31:0] _GEN_503;
  wire [31:0] _GEN_504;
  wire [31:0] _GEN_505;
  wire [31:0] _GEN_506;
  wire [31:0] _GEN_507;
  wire [31:0] _GEN_508;
  wire [31:0] _GEN_509;
  wire [31:0] _GEN_510;
  wire [31:0] _GEN_511;
  wire [31:0] _GEN_512;
  wire [31:0] _GEN_513;
  wire [31:0] _GEN_514;
  wire [31:0] _GEN_515;
  wire [31:0] _GEN_516;
  wire [31:0] _GEN_517;
  wire [31:0] _GEN_518;
  wire [31:0] _GEN_519;
  wire [31:0] _GEN_520;
  wire [31:0] _GEN_521;
  wire [31:0] _GEN_522;
  wire [31:0] _GEN_523;
  wire [31:0] _GEN_524;
  wire [31:0] _GEN_525;
  wire [31:0] _GEN_526;
  wire [31:0] _GEN_527;
  wire [31:0] _GEN_528;
  wire [31:0] _GEN_529;
  wire [31:0] _GEN_530;
  wire [31:0] _GEN_531;
  wire [31:0] _GEN_532;
  wire [31:0] _GEN_533;
  wire [31:0] _GEN_534;
  wire [31:0] _GEN_535;
  wire [31:0] _GEN_536;
  wire [31:0] _GEN_537;
  wire [31:0] _GEN_538;
  wire [31:0] _GEN_539;
  wire [31:0] _GEN_540;
  wire [31:0] _GEN_541;
  wire [31:0] _GEN_542;
  wire [31:0] _GEN_543;
  wire [31:0] _GEN_544;
  wire [31:0] _GEN_545;
  wire [31:0] _GEN_546;
  wire [31:0] _GEN_547;
  wire [31:0] _GEN_548;
  wire [31:0] _GEN_549;
  wire [31:0] _GEN_550;
  wire [31:0] _GEN_551;
  wire [31:0] _GEN_552;
  wire [31:0] _GEN_553;
  wire [31:0] _GEN_554;
  wire [31:0] _GEN_555;
  wire [31:0] _GEN_556;
  wire [31:0] _GEN_557;
  wire [31:0] _GEN_558;
  wire [31:0] _GEN_559;
  wire [31:0] _GEN_560;
  wire [31:0] _GEN_561;
  wire [31:0] _GEN_562;
  wire [31:0] _GEN_563;
  wire [31:0] _GEN_564;
  wire [31:0] _GEN_565;
  wire [31:0] _GEN_566;
  wire [31:0] _GEN_567;
  wire [31:0] _GEN_568;
  wire [31:0] _GEN_569;
  wire [31:0] _GEN_570;
  wire [31:0] _GEN_571;
  wire [31:0] _GEN_572;
  wire [31:0] _GEN_573;
  wire [31:0] _GEN_574;
  wire [31:0] _GEN_575;
  wire [31:0] _GEN_576;
  wire [31:0] _GEN_577;
  wire [31:0] _GEN_578;
  wire [31:0] _GEN_579;
  wire [31:0] _GEN_580;
  wire [31:0] _GEN_581;
  wire [31:0] _GEN_582;
  wire [31:0] _GEN_583;
  wire [31:0] _GEN_584;
  wire [31:0] _GEN_585;
  wire [31:0] _GEN_586;
  wire [31:0] _GEN_587;
  wire [31:0] _GEN_588;
  wire [31:0] _GEN_589;
  wire [31:0] _GEN_590;
  wire [31:0] _GEN_591;
  wire [31:0] _GEN_592;
  wire [31:0] _GEN_593;
  wire [31:0] _GEN_594;
  wire [31:0] _GEN_595;
  wire [31:0] _GEN_596;
  wire [31:0] _GEN_597;
  wire [31:0] _GEN_598;
  wire [31:0] _GEN_599;
  wire [31:0] _GEN_600;
  wire [31:0] _GEN_601;
  wire [31:0] _GEN_602;
  wire [31:0] _GEN_603;
  wire [31:0] _GEN_604;
  wire [31:0] _GEN_605;
  wire [31:0] _GEN_606;
  wire [31:0] _GEN_607;
  wire [31:0] _GEN_608;
  wire [31:0] _GEN_609;
  wire [31:0] _GEN_610;
  wire [31:0] _GEN_611;
  wire [31:0] _GEN_612;
  wire [31:0] _GEN_613;
  wire [31:0] _GEN_614;
  wire [31:0] _GEN_615;
  wire [31:0] _GEN_616;
  wire [31:0] _GEN_617;
  wire [31:0] _GEN_618;
  wire [31:0] _GEN_619;
  wire [31:0] _GEN_620;
  wire [31:0] _GEN_621;
  wire [31:0] _GEN_622;
  wire [31:0] _GEN_623;
  wire [31:0] _GEN_624;
  wire [31:0] _GEN_625;
  wire [31:0] _GEN_626;
  wire [31:0] _GEN_627;
  wire [31:0] _GEN_628;
  wire [31:0] _GEN_629;
  wire [31:0] _GEN_630;
  wire [31:0] _GEN_631;
  wire [31:0] _GEN_632;
  wire [31:0] _GEN_633;
  wire [31:0] _GEN_634;
  wire [31:0] _GEN_635;
  wire [31:0] _GEN_636;
  wire [31:0] _GEN_637;
  wire [31:0] _GEN_638;
  wire [31:0] _GEN_639;
  wire [31:0] _GEN_640;
  wire [31:0] _GEN_641;
  wire [31:0] _GEN_642;
  wire [31:0] _GEN_643;
  wire [31:0] _GEN_644;
  wire [31:0] _GEN_645;
  wire [31:0] _GEN_646;
  wire [31:0] _GEN_647;
  wire [31:0] _GEN_648;
  wire [31:0] _GEN_649;
  wire [31:0] _GEN_650;
  wire [31:0] _GEN_651;
  wire [31:0] _GEN_652;
  wire [31:0] _GEN_653;
  wire [31:0] _GEN_654;
  wire [31:0] _GEN_655;
  wire [31:0] _GEN_656;
  wire [31:0] _GEN_657;
  wire [31:0] _GEN_658;
  wire [31:0] _GEN_659;
  wire [31:0] _GEN_660;
  wire [31:0] _GEN_661;
  wire [31:0] _GEN_662;
  wire [31:0] _GEN_663;
  wire [31:0] _GEN_664;
  wire [31:0] _GEN_665;
  wire [31:0] _GEN_666;
  wire [31:0] _GEN_667;
  wire [31:0] _GEN_668;
  wire [31:0] _GEN_669;
  wire [31:0] _GEN_670;
  wire [31:0] _GEN_671;
  wire [31:0] _GEN_672;
  wire [31:0] _GEN_673;
  wire [31:0] _GEN_674;
  wire [31:0] _GEN_675;
  wire [31:0] _GEN_676;
  wire [31:0] _GEN_677;
  wire [31:0] _GEN_678;
  wire [31:0] _GEN_679;
  wire [31:0] _GEN_680;
  wire [31:0] _GEN_681;
  wire [31:0] _GEN_682;
  wire [31:0] _GEN_683;
  wire [31:0] _GEN_684;
  wire [31:0] _GEN_685;
  wire [31:0] _GEN_686;
  wire [31:0] _GEN_687;
  wire [31:0] _GEN_688;
  wire [31:0] _GEN_689;
  wire [31:0] _GEN_690;
  wire [31:0] _GEN_691;
  wire [31:0] _GEN_692;
  wire [31:0] _GEN_693;
  wire [31:0] _GEN_694;
  wire [31:0] _GEN_695;
  wire [31:0] _GEN_696;
  wire [31:0] _GEN_697;
  wire [31:0] _GEN_698;
  wire [31:0] _GEN_699;
  wire [31:0] _GEN_700;
  wire [31:0] _GEN_701;
  wire [31:0] _GEN_702;
  wire [31:0] _GEN_703;
  wire [31:0] _GEN_704;
  wire [31:0] _GEN_705;
  wire [31:0] _GEN_706;
  wire [31:0] _GEN_707;
  wire [31:0] _GEN_708;
  wire [31:0] _GEN_709;
  wire [31:0] _GEN_710;
  wire [31:0] _GEN_711;
  wire [31:0] _GEN_712;
  wire [31:0] _GEN_713;
  wire [31:0] _GEN_714;
  wire [31:0] _GEN_715;
  wire [31:0] _GEN_716;
  wire [31:0] _GEN_717;
  wire [31:0] _GEN_718;
  wire [31:0] _GEN_719;
  wire [31:0] _GEN_720;
  wire [31:0] _GEN_721;
  wire [31:0] _GEN_722;
  wire [31:0] _GEN_723;
  wire [31:0] _GEN_724;
  wire [31:0] _GEN_725;
  wire [31:0] _GEN_726;
  wire [31:0] _GEN_727;
  wire [31:0] _GEN_728;
  wire [31:0] _GEN_729;
  wire [31:0] _GEN_730;
  wire [31:0] _GEN_731;
  wire [31:0] _GEN_732;
  wire [31:0] _GEN_733;
  wire [31:0] _GEN_734;
  wire [31:0] _GEN_735;
  wire [31:0] _GEN_736;
  wire [31:0] _GEN_737;
  wire [31:0] _GEN_738;
  wire [31:0] _GEN_739;
  wire [31:0] _GEN_740;
  wire [31:0] _GEN_741;
  wire [31:0] _GEN_742;
  wire [31:0] _GEN_743;
  wire [31:0] _GEN_744;
  wire [31:0] _GEN_745;
  wire [31:0] _GEN_746;
  wire [31:0] _GEN_747;
  wire [31:0] _GEN_748;
  wire [31:0] _GEN_749;
  wire [31:0] _GEN_750;
  wire [31:0] _GEN_751;
  wire [31:0] _GEN_752;
  wire [31:0] _GEN_753;
  wire [31:0] _GEN_754;
  wire [31:0] _GEN_755;
  wire [31:0] _GEN_756;
  wire [31:0] _GEN_757;
  wire [31:0] _GEN_758;
  wire [31:0] _GEN_759;
  wire [31:0] _GEN_760;
  wire [31:0] _GEN_761;
  wire [31:0] _GEN_762;
  wire [31:0] _GEN_763;
  wire [31:0] _GEN_764;
  wire [31:0] _GEN_765;
  wire [31:0] _GEN_766;
  wire [31:0] _GEN_767;
  wire [31:0] _GEN_768;
  wire [31:0] _GEN_769;
  wire [31:0] _GEN_770;
  wire [31:0] _GEN_771;
  wire [31:0] _GEN_772;
  wire [31:0] _GEN_773;
  wire [31:0] _GEN_774;
  wire [31:0] _GEN_775;
  wire [31:0] _GEN_776;
  wire [31:0] _GEN_777;
  wire [31:0] _GEN_778;
  wire [31:0] _GEN_779;
  wire [31:0] _GEN_780;
  wire [31:0] _GEN_781;
  wire [31:0] _GEN_782;
  wire [31:0] _GEN_783;
  wire [31:0] _GEN_784;
  wire [31:0] _GEN_785;
  wire [31:0] _GEN_786;
  wire [31:0] _GEN_787;
  wire [31:0] _GEN_788;
  wire [31:0] _GEN_789;
  wire [31:0] _GEN_790;
  wire [31:0] _GEN_791;
  wire [31:0] _GEN_792;
  wire [31:0] _GEN_793;
  wire [31:0] _GEN_794;
  wire [31:0] _GEN_795;
  wire [31:0] _GEN_796;
  wire [31:0] _GEN_797;
  wire [31:0] _GEN_798;
  wire [31:0] _GEN_799;
  wire [31:0] _GEN_800;
  wire [31:0] _GEN_801;
  wire [31:0] _GEN_802;
  wire [31:0] _GEN_803;
  wire [31:0] _GEN_804;
  wire [31:0] _GEN_805;
  wire [31:0] _GEN_806;
  wire [31:0] _GEN_807;
  wire [31:0] _GEN_808;
  wire [31:0] _GEN_809;
  wire [31:0] _GEN_810;
  wire [31:0] _GEN_811;
  wire [31:0] _GEN_812;
  wire [31:0] _GEN_813;
  wire [31:0] _GEN_814;
  wire [31:0] _GEN_815;
  wire [31:0] _GEN_816;
  wire [31:0] _GEN_817;
  wire [31:0] _GEN_818;
  wire [31:0] _GEN_819;
  wire [31:0] _GEN_820;
  wire [31:0] _GEN_821;
  wire [31:0] _GEN_822;
  wire [31:0] _GEN_823;
  wire [31:0] _GEN_824;
  wire [31:0] _GEN_825;
  wire [31:0] _GEN_826;
  wire [31:0] _GEN_827;
  wire [31:0] _GEN_828;
  wire [31:0] _GEN_829;
  wire [31:0] _GEN_830;
  wire [31:0] _GEN_831;
  wire [31:0] _GEN_832;
  wire [31:0] _GEN_833;
  wire [31:0] _GEN_834;
  wire [31:0] _GEN_835;
  wire [31:0] _GEN_836;
  wire [31:0] _GEN_837;
  wire [31:0] _GEN_838;
  wire [31:0] _GEN_839;
  wire [31:0] _GEN_840;
  wire [31:0] _GEN_841;
  wire [31:0] _GEN_842;
  wire [31:0] _GEN_843;
  wire [31:0] _GEN_844;
  wire [31:0] _GEN_845;
  wire [31:0] _GEN_846;
  wire [31:0] _GEN_847;
  wire [31:0] _GEN_848;
  wire [31:0] _GEN_849;
  wire [31:0] _GEN_850;
  wire [31:0] _GEN_851;
  wire [31:0] _GEN_852;
  wire [31:0] _GEN_853;
  wire [31:0] _GEN_854;
  wire [31:0] _GEN_855;
  wire [31:0] _GEN_856;
  wire [31:0] _GEN_857;
  wire [31:0] _GEN_858;
  wire [31:0] _GEN_859;
  wire [31:0] _GEN_860;
  wire [31:0] _GEN_861;
  wire [31:0] _GEN_862;
  wire [31:0] _GEN_863;
  wire [31:0] _GEN_864;
  wire [31:0] _GEN_865;
  wire [31:0] _GEN_866;
  wire [31:0] _GEN_867;
  wire [31:0] _GEN_868;
  wire [31:0] _GEN_869;
  wire [31:0] _GEN_870;
  wire [31:0] _GEN_871;
  wire [31:0] _GEN_872;
  wire [31:0] _GEN_873;
  wire [31:0] _GEN_874;
  wire [31:0] _GEN_875;
  wire [31:0] _GEN_876;
  wire [31:0] _GEN_877;
  wire [31:0] _GEN_878;
  wire [31:0] _GEN_879;
  wire [31:0] _GEN_880;
  wire [31:0] _GEN_881;
  wire [31:0] _GEN_882;
  wire [31:0] _GEN_883;
  wire [31:0] _GEN_884;
  wire [31:0] _GEN_885;
  wire [31:0] _GEN_886;
  wire [31:0] _GEN_887;
  wire [31:0] _GEN_888;
  wire [31:0] _GEN_889;
  wire [31:0] _GEN_890;
  wire [31:0] _GEN_891;
  wire [31:0] _GEN_892;
  wire [31:0] _GEN_893;
  wire [31:0] _GEN_894;
  wire [31:0] _GEN_895;
  wire [31:0] _GEN_896;
  wire [31:0] _GEN_897;
  wire [31:0] _GEN_898;
  wire [31:0] _GEN_899;
  wire [31:0] _GEN_900;
  wire [31:0] _GEN_901;
  wire [31:0] _GEN_902;
  wire [31:0] _GEN_903;
  wire [31:0] _GEN_904;
  wire [31:0] _GEN_905;
  wire [31:0] _GEN_906;
  wire [31:0] _GEN_907;
  wire [31:0] _GEN_908;
  wire [31:0] _GEN_909;
  wire [31:0] _GEN_910;
  wire [31:0] _GEN_911;
  wire [31:0] _GEN_912;
  wire [31:0] _GEN_913;
  wire [31:0] _GEN_914;
  wire [31:0] _GEN_915;
  wire [31:0] _GEN_916;
  wire [31:0] _GEN_917;
  wire [31:0] _GEN_918;
  wire [31:0] _GEN_919;
  wire [31:0] _GEN_920;
  wire [31:0] _GEN_921;
  wire [31:0] _GEN_922;
  wire [31:0] _GEN_923;
  wire [31:0] _GEN_924;
  wire [31:0] _GEN_925;
  wire [31:0] _GEN_926;
  wire [31:0] _GEN_927;
  wire [31:0] _GEN_928;
  wire [31:0] _GEN_929;
  wire [31:0] _GEN_930;
  wire [31:0] _GEN_931;
  wire [31:0] _GEN_932;
  wire [31:0] _GEN_933;
  wire [31:0] _GEN_934;
  wire [31:0] _GEN_935;
  wire [31:0] _GEN_936;
  wire [31:0] _GEN_937;
  wire [31:0] _GEN_938;
  wire [31:0] _GEN_939;
  wire [31:0] _GEN_940;
  wire [31:0] _GEN_941;
  wire [31:0] _GEN_942;
  wire [31:0] _GEN_943;
  wire [31:0] _GEN_944;
  wire [31:0] _GEN_945;
  wire [31:0] _GEN_946;
  wire [31:0] _GEN_947;
  wire [31:0] _GEN_948;
  wire [31:0] _GEN_949;
  wire [31:0] _GEN_950;
  wire [31:0] _GEN_951;
  wire [31:0] _GEN_952;
  wire [31:0] _GEN_953;
  wire [31:0] _GEN_954;
  wire [31:0] _GEN_955;
  wire [31:0] _GEN_956;
  wire [31:0] _GEN_957;
  wire [31:0] _GEN_958;
  wire [31:0] _GEN_959;
  wire [31:0] _GEN_960;
  wire [31:0] _GEN_961;
  wire [31:0] _GEN_962;
  wire [31:0] _GEN_963;
  wire [31:0] _GEN_964;
  wire [31:0] _GEN_965;
  wire [31:0] _GEN_966;
  wire [31:0] _GEN_967;
  wire [31:0] _GEN_968;
  wire [31:0] _GEN_969;
  wire [31:0] _GEN_970;
  wire [31:0] _GEN_971;
  wire [31:0] _GEN_972;
  wire [31:0] _GEN_973;
  wire [31:0] _GEN_974;
  wire [31:0] _GEN_975;
  wire [31:0] _GEN_976;
  wire [31:0] _GEN_977;
  wire [31:0] _GEN_978;
  wire [31:0] _GEN_979;
  wire [31:0] _GEN_980;
  wire [31:0] _GEN_981;
  wire [31:0] _GEN_982;
  wire [31:0] _GEN_983;
  wire [31:0] _GEN_984;
  wire [31:0] _GEN_985;
  wire [31:0] _GEN_986;
  wire [31:0] _GEN_987;
  wire [31:0] _GEN_988;
  wire [31:0] _GEN_989;
  wire [31:0] _GEN_990;
  wire [31:0] _GEN_991;
  wire [31:0] _GEN_992;
  wire [31:0] _GEN_993;
  wire [31:0] _GEN_994;
  wire [31:0] _GEN_995;
  wire [31:0] _GEN_996;
  wire [31:0] _GEN_997;
  wire [31:0] _GEN_998;
  wire [31:0] _GEN_999;
  wire [31:0] _GEN_1000;
  wire [31:0] _GEN_1001;
  wire [31:0] _GEN_1002;
  wire [31:0] _GEN_1003;
  wire [31:0] _GEN_1004;
  wire [31:0] _GEN_1005;
  wire [31:0] _GEN_1006;
  wire [31:0] _GEN_1007;
  wire [31:0] _GEN_1008;
  wire [31:0] _GEN_1009;
  wire [31:0] _GEN_1010;
  wire [31:0] _GEN_1011;
  wire [31:0] _GEN_1012;
  wire [31:0] _GEN_1013;
  wire [31:0] _GEN_1014;
  wire [31:0] _GEN_1015;
  wire [31:0] _GEN_1016;
  wire [31:0] _GEN_1017;
  wire [31:0] _GEN_1018;
  wire [31:0] _GEN_1019;
  wire [31:0] _GEN_1020;
  wire [31:0] _GEN_1021;
  wire [31:0] _GEN_1022;
  wire [31:0] _GEN_1023;
  wire [31:0] _T_2116;
  assign io_in_0_a_ready = io_in_0_d_ready;
  assign io_in_0_d_valid = io_in_0_a_valid;
  assign io_in_0_d_bits_opcode = 3'h1;
  assign io_in_0_d_bits_param = 2'h0;
  assign io_in_0_d_bits_size = io_in_0_a_bits_size;
  assign io_in_0_d_bits_source = io_in_0_a_bits_source;
  assign io_in_0_d_bits_sink = 1'h0;
  assign io_in_0_d_bits_data = _T_2116;
  assign io_in_0_d_bits_error = 1'h0;
  assign index = io_in_0_a_bits_address[11:2];
  assign high = io_in_0_a_bits_address[15:12];
  assign _T_2113 = high != 4'h0;
  assign _GEN_1 = 10'h1 == index ? 32'h1f41413 : 32'h10041b;
  assign _GEN_2 = 10'h2 == index ? 32'hf1402573 : _GEN_1;
  assign _GEN_3 = 10'h3 == index ? 32'h597 : _GEN_2;
  assign _GEN_4 = 10'h4 == index ? 32'h7458593 : _GEN_3;
  assign _GEN_5 = 10'h5 == index ? 32'h8402 : _GEN_4;
  assign _GEN_6 = 10'h6 == index ? 32'h0 : _GEN_5;
  assign _GEN_7 = 10'h7 == index ? 32'h0 : _GEN_6;
  assign _GEN_8 = 10'h8 == index ? 32'h0 : _GEN_7;
  assign _GEN_9 = 10'h9 == index ? 32'h0 : _GEN_8;
  assign _GEN_10 = 10'ha == index ? 32'h0 : _GEN_9;
  assign _GEN_11 = 10'hb == index ? 32'h0 : _GEN_10;
  assign _GEN_12 = 10'hc == index ? 32'h0 : _GEN_11;
  assign _GEN_13 = 10'hd == index ? 32'h0 : _GEN_12;
  assign _GEN_14 = 10'he == index ? 32'h0 : _GEN_13;
  assign _GEN_15 = 10'hf == index ? 32'h0 : _GEN_14;
  assign _GEN_16 = 10'h10 == index ? 32'hf1402573 : _GEN_15;
  assign _GEN_17 = 10'h11 == index ? 32'h597 : _GEN_16;
  assign _GEN_18 = 10'h12 == index ? 32'h3c58593 : _GEN_17;
  assign _GEN_19 = 10'h13 == index ? 32'h10500073 : _GEN_18;
  assign _GEN_20 = 10'h14 == index ? 32'hbff5 : _GEN_19;
  assign _GEN_21 = 10'h15 == index ? 32'h0 : _GEN_20;
  assign _GEN_22 = 10'h16 == index ? 32'h0 : _GEN_21;
  assign _GEN_23 = 10'h17 == index ? 32'h0 : _GEN_22;
  assign _GEN_24 = 10'h18 == index ? 32'h0 : _GEN_23;
  assign _GEN_25 = 10'h19 == index ? 32'h0 : _GEN_24;
  assign _GEN_26 = 10'h1a == index ? 32'h0 : _GEN_25;
  assign _GEN_27 = 10'h1b == index ? 32'h0 : _GEN_26;
  assign _GEN_28 = 10'h1c == index ? 32'h0 : _GEN_27;
  assign _GEN_29 = 10'h1d == index ? 32'h0 : _GEN_28;
  assign _GEN_30 = 10'h1e == index ? 32'h0 : _GEN_29;
  assign _GEN_31 = 10'h1f == index ? 32'h0 : _GEN_30;
  assign _GEN_32 = 10'h20 == index ? 32'hedfe0dd0 : _GEN_31;
  assign _GEN_33 = 10'h21 == index ? 32'hdd070000 : _GEN_32;
  assign _GEN_34 = 10'h22 == index ? 32'h38000000 : _GEN_33;
  assign _GEN_35 = 10'h23 == index ? 32'h90060000 : _GEN_34;
  assign _GEN_36 = 10'h24 == index ? 32'h28000000 : _GEN_35;
  assign _GEN_37 = 10'h25 == index ? 32'h11000000 : _GEN_36;
  assign _GEN_38 = 10'h26 == index ? 32'h10000000 : _GEN_37;
  assign _GEN_39 = 10'h27 == index ? 32'h0 : _GEN_38;
  assign _GEN_40 = 10'h28 == index ? 32'h4d010000 : _GEN_39;
  assign _GEN_41 = 10'h29 == index ? 32'h58060000 : _GEN_40;
  assign _GEN_42 = 10'h2a == index ? 32'h0 : _GEN_41;
  assign _GEN_43 = 10'h2b == index ? 32'h0 : _GEN_42;
  assign _GEN_44 = 10'h2c == index ? 32'h0 : _GEN_43;
  assign _GEN_45 = 10'h2d == index ? 32'h0 : _GEN_44;
  assign _GEN_46 = 10'h2e == index ? 32'h1000000 : _GEN_45;
  assign _GEN_47 = 10'h2f == index ? 32'h0 : _GEN_46;
  assign _GEN_48 = 10'h30 == index ? 32'h3000000 : _GEN_47;
  assign _GEN_49 = 10'h31 == index ? 32'h4000000 : _GEN_48;
  assign _GEN_50 = 10'h32 == index ? 32'h0 : _GEN_49;
  assign _GEN_51 = 10'h33 == index ? 32'h1000000 : _GEN_50;
  assign _GEN_52 = 10'h34 == index ? 32'h3000000 : _GEN_51;
  assign _GEN_53 = 10'h35 == index ? 32'h4000000 : _GEN_52;
  assign _GEN_54 = 10'h36 == index ? 32'hf000000 : _GEN_53;
  assign _GEN_55 = 10'h37 == index ? 32'h1000000 : _GEN_54;
  assign _GEN_56 = 10'h38 == index ? 32'h3000000 : _GEN_55;
  assign _GEN_57 = 10'h39 == index ? 32'h21000000 : _GEN_56;
  assign _GEN_58 = 10'h3a == index ? 32'h1b000000 : _GEN_57;
  assign _GEN_59 = 10'h3b == index ? 32'h65657266 : _GEN_58;
  assign _GEN_60 = 10'h3c == index ? 32'h70696863 : _GEN_59;
  assign _GEN_61 = 10'h3d == index ? 32'h6f722c73 : _GEN_60;
  assign _GEN_62 = 10'h3e == index ? 32'h74656b63 : _GEN_61;
  assign _GEN_63 = 10'h3f == index ? 32'h70696863 : _GEN_62;
  assign _GEN_64 = 10'h40 == index ? 32'h6b6e752d : _GEN_63;
  assign _GEN_65 = 10'h41 == index ? 32'h6e776f6e : _GEN_64;
  assign _GEN_66 = 10'h42 == index ? 32'h7665642d : _GEN_65;
  assign _GEN_67 = 10'h43 == index ? 32'h0 : _GEN_66;
  assign _GEN_68 = 10'h44 == index ? 32'h3000000 : _GEN_67;
  assign _GEN_69 = 10'h45 == index ? 32'h1d000000 : _GEN_68;
  assign _GEN_70 = 10'h46 == index ? 32'h26000000 : _GEN_69;
  assign _GEN_71 = 10'h47 == index ? 32'h65657266 : _GEN_70;
  assign _GEN_72 = 10'h48 == index ? 32'h70696863 : _GEN_71;
  assign _GEN_73 = 10'h49 == index ? 32'h6f722c73 : _GEN_72;
  assign _GEN_74 = 10'h4a == index ? 32'h74656b63 : _GEN_73;
  assign _GEN_75 = 10'h4b == index ? 32'h70696863 : _GEN_74;
  assign _GEN_76 = 10'h4c == index ? 32'h6b6e752d : _GEN_75;
  assign _GEN_77 = 10'h4d == index ? 32'h6e776f6e : _GEN_76;
  assign _GEN_78 = 10'h4e == index ? 32'h0 : _GEN_77;
  assign _GEN_79 = 10'h4f == index ? 32'h1000000 : _GEN_78;
  assign _GEN_80 = 10'h50 == index ? 32'h73757063 : _GEN_79;
  assign _GEN_81 = 10'h51 == index ? 32'h0 : _GEN_80;
  assign _GEN_82 = 10'h52 == index ? 32'h3000000 : _GEN_81;
  assign _GEN_83 = 10'h53 == index ? 32'h4000000 : _GEN_82;
  assign _GEN_84 = 10'h54 == index ? 32'h0 : _GEN_83;
  assign _GEN_85 = 10'h55 == index ? 32'h1000000 : _GEN_84;
  assign _GEN_86 = 10'h56 == index ? 32'h3000000 : _GEN_85;
  assign _GEN_87 = 10'h57 == index ? 32'h4000000 : _GEN_86;
  assign _GEN_88 = 10'h58 == index ? 32'hf000000 : _GEN_87;
  assign _GEN_89 = 10'h59 == index ? 32'h0 : _GEN_88;
  assign _GEN_90 = 10'h5a == index ? 32'h3000000 : _GEN_89;
  assign _GEN_91 = 10'h5b == index ? 32'h4000000 : _GEN_90;
  assign _GEN_92 = 10'h5c == index ? 32'h2c000000 : _GEN_91;
  assign _GEN_93 = 10'h5d == index ? 32'h40420f00 : _GEN_92;
  assign _GEN_94 = 10'h5e == index ? 32'h1000000 : _GEN_93;
  assign _GEN_95 = 10'h5f == index ? 32'h40757063 : _GEN_94;
  assign _GEN_96 = 10'h60 == index ? 32'h30 : _GEN_95;
  assign _GEN_97 = 10'h61 == index ? 32'h3000000 : _GEN_96;
  assign _GEN_98 = 10'h62 == index ? 32'h4000000 : _GEN_97;
  assign _GEN_99 = 10'h63 == index ? 32'h3f000000 : _GEN_98;
  assign _GEN_100 = 10'h64 == index ? 32'h0 : _GEN_99;
  assign _GEN_101 = 10'h65 == index ? 32'h3000000 : _GEN_100;
  assign _GEN_102 = 10'h66 == index ? 32'h15000000 : _GEN_101;
  assign _GEN_103 = 10'h67 == index ? 32'h1b000000 : _GEN_102;
  assign _GEN_104 = 10'h68 == index ? 32'h69666973 : _GEN_103;
  assign _GEN_105 = 10'h69 == index ? 32'h722c6576 : _GEN_104;
  assign _GEN_106 = 10'h6a == index ? 32'h656b636f : _GEN_105;
  assign _GEN_107 = 10'h6b == index ? 32'h72003074 : _GEN_106;
  assign _GEN_108 = 10'h6c == index ? 32'h76637369 : _GEN_107;
  assign _GEN_109 = 10'h6d == index ? 32'h0 : _GEN_108;
  assign _GEN_110 = 10'h6e == index ? 32'h3000000 : _GEN_109;
  assign _GEN_111 = 10'h6f == index ? 32'h4000000 : _GEN_110;
  assign _GEN_112 = 10'h70 == index ? 32'h4f000000 : _GEN_111;
  assign _GEN_113 = 10'h71 == index ? 32'h757063 : _GEN_112;
  assign _GEN_114 = 10'h72 == index ? 32'h3000000 : _GEN_113;
  assign _GEN_115 = 10'h73 == index ? 32'h4000000 : _GEN_114;
  assign _GEN_116 = 10'h74 == index ? 32'h5b000000 : _GEN_115;
  assign _GEN_117 = 10'h75 == index ? 32'h40000000 : _GEN_116;
  assign _GEN_118 = 10'h76 == index ? 32'h3000000 : _GEN_117;
  assign _GEN_119 = 10'h77 == index ? 32'h4000000 : _GEN_118;
  assign _GEN_120 = 10'h78 == index ? 32'h6e000000 : _GEN_119;
  assign _GEN_121 = 10'h79 == index ? 32'h40000000 : _GEN_120;
  assign _GEN_122 = 10'h7a == index ? 32'h3000000 : _GEN_121;
  assign _GEN_123 = 10'h7b == index ? 32'h4000000 : _GEN_122;
  assign _GEN_124 = 10'h7c == index ? 32'h7b000000 : _GEN_123;
  assign _GEN_125 = 10'h7d == index ? 32'h100000 : _GEN_124;
  assign _GEN_126 = 10'h7e == index ? 32'h3000000 : _GEN_125;
  assign _GEN_127 = 10'h7f == index ? 32'h4000000 : _GEN_126;
  assign _GEN_128 = 10'h80 == index ? 32'h88000000 : _GEN_127;
  assign _GEN_129 = 10'h81 == index ? 32'h1000000 : _GEN_128;
  assign _GEN_130 = 10'h82 == index ? 32'h3000000 : _GEN_129;
  assign _GEN_131 = 10'h83 == index ? 32'h4000000 : _GEN_130;
  assign _GEN_132 = 10'h84 == index ? 32'h99000000 : _GEN_131;
  assign _GEN_133 = 10'h85 == index ? 32'h0 : _GEN_132;
  assign _GEN_134 = 10'h86 == index ? 32'h3000000 : _GEN_133;
  assign _GEN_135 = 10'h87 == index ? 32'h9000000 : _GEN_134;
  assign _GEN_136 = 10'h88 == index ? 32'h9d000000 : _GEN_135;
  assign _GEN_137 = 10'h89 == index ? 32'h32337672 : _GEN_136;
  assign _GEN_138 = 10'h8a == index ? 32'h63616d69 : _GEN_137;
  assign _GEN_139 = 10'h8b == index ? 32'h0 : _GEN_138;
  assign _GEN_140 = 10'h8c == index ? 32'h3000000 : _GEN_139;
  assign _GEN_141 = 10'h8d == index ? 32'h4000000 : _GEN_140;
  assign _GEN_142 = 10'h8e == index ? 32'ha7000000 : _GEN_141;
  assign _GEN_143 = 10'h8f == index ? 32'h2000000 : _GEN_142;
  assign _GEN_144 = 10'h90 == index ? 32'h3000000 : _GEN_143;
  assign _GEN_145 = 10'h91 == index ? 32'h5000000 : _GEN_144;
  assign _GEN_146 = 10'h92 == index ? 32'hb3000000 : _GEN_145;
  assign _GEN_147 = 10'h93 == index ? 32'h79616b6f : _GEN_146;
  assign _GEN_148 = 10'h94 == index ? 32'h0 : _GEN_147;
  assign _GEN_149 = 10'h95 == index ? 32'h1000000 : _GEN_148;
  assign _GEN_150 = 10'h96 == index ? 32'h65746e69 : _GEN_149;
  assign _GEN_151 = 10'h97 == index ? 32'h70757272 : _GEN_150;
  assign _GEN_152 = 10'h98 == index ? 32'h6f632d74 : _GEN_151;
  assign _GEN_153 = 10'h99 == index ? 32'h6f72746e : _GEN_152;
  assign _GEN_154 = 10'h9a == index ? 32'h72656c6c : _GEN_153;
  assign _GEN_155 = 10'h9b == index ? 32'h0 : _GEN_154;
  assign _GEN_156 = 10'h9c == index ? 32'h3000000 : _GEN_155;
  assign _GEN_157 = 10'h9d == index ? 32'h4000000 : _GEN_156;
  assign _GEN_158 = 10'h9e == index ? 32'hba000000 : _GEN_157;
  assign _GEN_159 = 10'h9f == index ? 32'h1000000 : _GEN_158;
  assign _GEN_160 = 10'ha0 == index ? 32'h3000000 : _GEN_159;
  assign _GEN_161 = 10'ha1 == index ? 32'hf000000 : _GEN_160;
  assign _GEN_162 = 10'ha2 == index ? 32'h1b000000 : _GEN_161;
  assign _GEN_163 = 10'ha3 == index ? 32'h63736972 : _GEN_162;
  assign _GEN_164 = 10'ha4 == index ? 32'h70632c76 : _GEN_163;
  assign _GEN_165 = 10'ha5 == index ? 32'h6e692d75 : _GEN_164;
  assign _GEN_166 = 10'ha6 == index ? 32'h6374 : _GEN_165;
  assign _GEN_167 = 10'ha7 == index ? 32'h3000000 : _GEN_166;
  assign _GEN_168 = 10'ha8 == index ? 32'h0 : _GEN_167;
  assign _GEN_169 = 10'ha9 == index ? 32'hcb000000 : _GEN_168;
  assign _GEN_170 = 10'haa == index ? 32'h3000000 : _GEN_169;
  assign _GEN_171 = 10'hab == index ? 32'h4000000 : _GEN_170;
  assign _GEN_172 = 10'hac == index ? 32'he0000000 : _GEN_171;
  assign _GEN_173 = 10'had == index ? 32'h3000000 : _GEN_172;
  assign _GEN_174 = 10'hae == index ? 32'h3000000 : _GEN_173;
  assign _GEN_175 = 10'haf == index ? 32'h4000000 : _GEN_174;
  assign _GEN_176 = 10'hb0 == index ? 32'he6000000 : _GEN_175;
  assign _GEN_177 = 10'hb1 == index ? 32'h3000000 : _GEN_176;
  assign _GEN_178 = 10'hb2 == index ? 32'h2000000 : _GEN_177;
  assign _GEN_179 = 10'hb3 == index ? 32'h2000000 : _GEN_178;
  assign _GEN_180 = 10'hb4 == index ? 32'h2000000 : _GEN_179;
  assign _GEN_181 = 10'hb5 == index ? 32'h1000000 : _GEN_180;
  assign _GEN_182 = 10'hb6 == index ? 32'h636f73 : _GEN_181;
  assign _GEN_183 = 10'hb7 == index ? 32'h3000000 : _GEN_182;
  assign _GEN_184 = 10'hb8 == index ? 32'h4000000 : _GEN_183;
  assign _GEN_185 = 10'hb9 == index ? 32'h0 : _GEN_184;
  assign _GEN_186 = 10'hba == index ? 32'h1000000 : _GEN_185;
  assign _GEN_187 = 10'hbb == index ? 32'h3000000 : _GEN_186;
  assign _GEN_188 = 10'hbc == index ? 32'h4000000 : _GEN_187;
  assign _GEN_189 = 10'hbd == index ? 32'hf000000 : _GEN_188;
  assign _GEN_190 = 10'hbe == index ? 32'h1000000 : _GEN_189;
  assign _GEN_191 = 10'hbf == index ? 32'h3000000 : _GEN_190;
  assign _GEN_192 = 10'hc0 == index ? 32'h2c000000 : _GEN_191;
  assign _GEN_193 = 10'hc1 == index ? 32'h1b000000 : _GEN_192;
  assign _GEN_194 = 10'hc2 == index ? 32'h65657266 : _GEN_193;
  assign _GEN_195 = 10'hc3 == index ? 32'h70696863 : _GEN_194;
  assign _GEN_196 = 10'hc4 == index ? 32'h6f722c73 : _GEN_195;
  assign _GEN_197 = 10'hc5 == index ? 32'h74656b63 : _GEN_196;
  assign _GEN_198 = 10'hc6 == index ? 32'h70696863 : _GEN_197;
  assign _GEN_199 = 10'hc7 == index ? 32'h6b6e752d : _GEN_198;
  assign _GEN_200 = 10'hc8 == index ? 32'h6e776f6e : _GEN_199;
  assign _GEN_201 = 10'hc9 == index ? 32'h636f732d : _GEN_200;
  assign _GEN_202 = 10'hca == index ? 32'h6d697300 : _GEN_201;
  assign _GEN_203 = 10'hcb == index ? 32'h2d656c70 : _GEN_202;
  assign _GEN_204 = 10'hcc == index ? 32'h737562 : _GEN_203;
  assign _GEN_205 = 10'hcd == index ? 32'h3000000 : _GEN_204;
  assign _GEN_206 = 10'hce == index ? 32'h0 : _GEN_205;
  assign _GEN_207 = 10'hcf == index ? 32'hee000000 : _GEN_206;
  assign _GEN_208 = 10'hd0 == index ? 32'h1000000 : _GEN_207;
  assign _GEN_209 = 10'hd1 == index ? 32'h6e696c63 : _GEN_208;
  assign _GEN_210 = 10'hd2 == index ? 32'h30324074 : _GEN_209;
  assign _GEN_211 = 10'hd3 == index ? 32'h30303030 : _GEN_210;
  assign _GEN_212 = 10'hd4 == index ? 32'h30 : _GEN_211;
  assign _GEN_213 = 10'hd5 == index ? 32'h3000000 : _GEN_212;
  assign _GEN_214 = 10'hd6 == index ? 32'hd000000 : _GEN_213;
  assign _GEN_215 = 10'hd7 == index ? 32'h1b000000 : _GEN_214;
  assign _GEN_216 = 10'hd8 == index ? 32'h63736972 : _GEN_215;
  assign _GEN_217 = 10'hd9 == index ? 32'h6c632c76 : _GEN_216;
  assign _GEN_218 = 10'hda == index ? 32'h30746e69 : _GEN_217;
  assign _GEN_219 = 10'hdb == index ? 32'h0 : _GEN_218;
  assign _GEN_220 = 10'hdc == index ? 32'h3000000 : _GEN_219;
  assign _GEN_221 = 10'hdd == index ? 32'h10000000 : _GEN_220;
  assign _GEN_222 = 10'hde == index ? 32'hf5000000 : _GEN_221;
  assign _GEN_223 = 10'hdf == index ? 32'h3000000 : _GEN_222;
  assign _GEN_224 = 10'he0 == index ? 32'h3000000 : _GEN_223;
  assign _GEN_225 = 10'he1 == index ? 32'h3000000 : _GEN_224;
  assign _GEN_226 = 10'he2 == index ? 32'h7000000 : _GEN_225;
  assign _GEN_227 = 10'he3 == index ? 32'h3000000 : _GEN_226;
  assign _GEN_228 = 10'he4 == index ? 32'h8000000 : _GEN_227;
  assign _GEN_229 = 10'he5 == index ? 32'h99000000 : _GEN_228;
  assign _GEN_230 = 10'he6 == index ? 32'h2 : _GEN_229;
  assign _GEN_231 = 10'he7 == index ? 32'h100 : _GEN_230;
  assign _GEN_232 = 10'he8 == index ? 32'h3000000 : _GEN_231;
  assign _GEN_233 = 10'he9 == index ? 32'h8000000 : _GEN_232;
  assign _GEN_234 = 10'hea == index ? 32'h9010000 : _GEN_233;
  assign _GEN_235 = 10'heb == index ? 32'h746e6f63 : _GEN_234;
  assign _GEN_236 = 10'hec == index ? 32'h6c6f72 : _GEN_235;
  assign _GEN_237 = 10'hed == index ? 32'h2000000 : _GEN_236;
  assign _GEN_238 = 10'hee == index ? 32'h1000000 : _GEN_237;
  assign _GEN_239 = 10'hef == index ? 32'h75626564 : _GEN_238;
  assign _GEN_240 = 10'hf0 == index ? 32'h6f632d67 : _GEN_239;
  assign _GEN_241 = 10'hf1 == index ? 32'h6f72746e : _GEN_240;
  assign _GEN_242 = 10'hf2 == index ? 32'h72656c6c : _GEN_241;
  assign _GEN_243 = 10'hf3 == index ? 32'h3040 : _GEN_242;
  assign _GEN_244 = 10'hf4 == index ? 32'h3000000 : _GEN_243;
  assign _GEN_245 = 10'hf5 == index ? 32'h21000000 : _GEN_244;
  assign _GEN_246 = 10'hf6 == index ? 32'h1b000000 : _GEN_245;
  assign _GEN_247 = 10'hf7 == index ? 32'h69666973 : _GEN_246;
  assign _GEN_248 = 10'hf8 == index ? 32'h642c6576 : _GEN_247;
  assign _GEN_249 = 10'hf9 == index ? 32'h67756265 : _GEN_248;
  assign _GEN_250 = 10'hfa == index ? 32'h3331302d : _GEN_249;
  assign _GEN_251 = 10'hfb == index ? 32'h73697200 : _GEN_250;
  assign _GEN_252 = 10'hfc == index ? 32'h642c7663 : _GEN_251;
  assign _GEN_253 = 10'hfd == index ? 32'h67756265 : _GEN_252;
  assign _GEN_254 = 10'hfe == index ? 32'h3331302d : _GEN_253;
  assign _GEN_255 = 10'hff == index ? 32'h0 : _GEN_254;
  assign _GEN_256 = 10'h100 == index ? 32'h3000000 : _GEN_255;
  assign _GEN_257 = 10'h101 == index ? 32'h8000000 : _GEN_256;
  assign _GEN_258 = 10'h102 == index ? 32'hf5000000 : _GEN_257;
  assign _GEN_259 = 10'h103 == index ? 32'h3000000 : _GEN_258;
  assign _GEN_260 = 10'h104 == index ? 32'hffff0000 : _GEN_259;
  assign _GEN_261 = 10'h105 == index ? 32'h3000000 : _GEN_260;
  assign _GEN_262 = 10'h106 == index ? 32'h8000000 : _GEN_261;
  assign _GEN_263 = 10'h107 == index ? 32'h99000000 : _GEN_262;
  assign _GEN_264 = 10'h108 == index ? 32'h0 : _GEN_263;
  assign _GEN_265 = 10'h109 == index ? 32'h100000 : _GEN_264;
  assign _GEN_266 = 10'h10a == index ? 32'h3000000 : _GEN_265;
  assign _GEN_267 = 10'h10b == index ? 32'h8000000 : _GEN_266;
  assign _GEN_268 = 10'h10c == index ? 32'h9010000 : _GEN_267;
  assign _GEN_269 = 10'h10d == index ? 32'h746e6f63 : _GEN_268;
  assign _GEN_270 = 10'h10e == index ? 32'h6c6f72 : _GEN_269;
  assign _GEN_271 = 10'h10f == index ? 32'h2000000 : _GEN_270;
  assign _GEN_272 = 10'h110 == index ? 32'h1000000 : _GEN_271;
  assign _GEN_273 = 10'h111 == index ? 32'h6d697464 : _GEN_272;
  assign _GEN_274 = 10'h112 == index ? 32'h30303840 : _GEN_273;
  assign _GEN_275 = 10'h113 == index ? 32'h30303030 : _GEN_274;
  assign _GEN_276 = 10'h114 == index ? 32'h30 : _GEN_275;
  assign _GEN_277 = 10'h115 == index ? 32'h3000000 : _GEN_276;
  assign _GEN_278 = 10'h116 == index ? 32'hd000000 : _GEN_277;
  assign _GEN_279 = 10'h117 == index ? 32'h1b000000 : _GEN_278;
  assign _GEN_280 = 10'h118 == index ? 32'h69666973 : _GEN_279;
  assign _GEN_281 = 10'h119 == index ? 32'h642c6576 : _GEN_280;
  assign _GEN_282 = 10'h11a == index ? 32'h306d6974 : _GEN_281;
  assign _GEN_283 = 10'h11b == index ? 32'h0 : _GEN_282;
  assign _GEN_284 = 10'h11c == index ? 32'h3000000 : _GEN_283;
  assign _GEN_285 = 10'h11d == index ? 32'h8000000 : _GEN_284;
  assign _GEN_286 = 10'h11e == index ? 32'h99000000 : _GEN_285;
  assign _GEN_287 = 10'h11f == index ? 32'h80 : _GEN_286;
  assign _GEN_288 = 10'h120 == index ? 32'h400000 : _GEN_287;
  assign _GEN_289 = 10'h121 == index ? 32'h3000000 : _GEN_288;
  assign _GEN_290 = 10'h122 == index ? 32'h4000000 : _GEN_289;
  assign _GEN_291 = 10'h123 == index ? 32'h9010000 : _GEN_290;
  assign _GEN_292 = 10'h124 == index ? 32'h6d656d : _GEN_291;
  assign _GEN_293 = 10'h125 == index ? 32'h3000000 : _GEN_292;
  assign _GEN_294 = 10'h126 == index ? 32'h4000000 : _GEN_293;
  assign _GEN_295 = 10'h127 == index ? 32'he0000000 : _GEN_294;
  assign _GEN_296 = 10'h128 == index ? 32'h2000000 : _GEN_295;
  assign _GEN_297 = 10'h129 == index ? 32'h3000000 : _GEN_296;
  assign _GEN_298 = 10'h12a == index ? 32'h4000000 : _GEN_297;
  assign _GEN_299 = 10'h12b == index ? 32'he6000000 : _GEN_298;
  assign _GEN_300 = 10'h12c == index ? 32'h2000000 : _GEN_299;
  assign _GEN_301 = 10'h12d == index ? 32'h2000000 : _GEN_300;
  assign _GEN_302 = 10'h12e == index ? 32'h1000000 : _GEN_301;
  assign _GEN_303 = 10'h12f == index ? 32'h6f727265 : _GEN_302;
  assign _GEN_304 = 10'h130 == index ? 32'h65642d72 : _GEN_303;
  assign _GEN_305 = 10'h131 == index ? 32'h65636976 : _GEN_304;
  assign _GEN_306 = 10'h132 == index ? 32'h30303340 : _GEN_305;
  assign _GEN_307 = 10'h133 == index ? 32'h30 : _GEN_306;
  assign _GEN_308 = 10'h134 == index ? 32'h3000000 : _GEN_307;
  assign _GEN_309 = 10'h135 == index ? 32'he000000 : _GEN_308;
  assign _GEN_310 = 10'h136 == index ? 32'h1b000000 : _GEN_309;
  assign _GEN_311 = 10'h137 == index ? 32'h69666973 : _GEN_310;
  assign _GEN_312 = 10'h138 == index ? 32'h652c6576 : _GEN_311;
  assign _GEN_313 = 10'h139 == index ? 32'h726f7272 : _GEN_312;
  assign _GEN_314 = 10'h13a == index ? 32'h30 : _GEN_313;
  assign _GEN_315 = 10'h13b == index ? 32'h3000000 : _GEN_314;
  assign _GEN_316 = 10'h13c == index ? 32'h8000000 : _GEN_315;
  assign _GEN_317 = 10'h13d == index ? 32'h99000000 : _GEN_316;
  assign _GEN_318 = 10'h13e == index ? 32'h300000 : _GEN_317;
  assign _GEN_319 = 10'h13f == index ? 32'h100000 : _GEN_318;
  assign _GEN_320 = 10'h140 == index ? 32'h3000000 : _GEN_319;
  assign _GEN_321 = 10'h141 == index ? 32'h4000000 : _GEN_320;
  assign _GEN_322 = 10'h142 == index ? 32'h9010000 : _GEN_321;
  assign _GEN_323 = 10'h143 == index ? 32'h6d656d : _GEN_322;
  assign _GEN_324 = 10'h144 == index ? 32'h3000000 : _GEN_323;
  assign _GEN_325 = 10'h145 == index ? 32'h4000000 : _GEN_324;
  assign _GEN_326 = 10'h146 == index ? 32'he0000000 : _GEN_325;
  assign _GEN_327 = 10'h147 == index ? 32'h1000000 : _GEN_326;
  assign _GEN_328 = 10'h148 == index ? 32'h3000000 : _GEN_327;
  assign _GEN_329 = 10'h149 == index ? 32'h4000000 : _GEN_328;
  assign _GEN_330 = 10'h14a == index ? 32'he6000000 : _GEN_329;
  assign _GEN_331 = 10'h14b == index ? 32'h1000000 : _GEN_330;
  assign _GEN_332 = 10'h14c == index ? 32'h2000000 : _GEN_331;
  assign _GEN_333 = 10'h14d == index ? 32'h1000000 : _GEN_332;
  assign _GEN_334 = 10'h14e == index ? 32'h65747865 : _GEN_333;
  assign _GEN_335 = 10'h14f == index ? 32'h6c616e72 : _GEN_334;
  assign _GEN_336 = 10'h150 == index ? 32'h746e692d : _GEN_335;
  assign _GEN_337 = 10'h151 == index ? 32'h75727265 : _GEN_336;
  assign _GEN_338 = 10'h152 == index ? 32'h737470 : _GEN_337;
  assign _GEN_339 = 10'h153 == index ? 32'h3000000 : _GEN_338;
  assign _GEN_340 = 10'h154 == index ? 32'h4000000 : _GEN_339;
  assign _GEN_341 = 10'h155 == index ? 32'h13010000 : _GEN_340;
  assign _GEN_342 = 10'h156 == index ? 32'h4000000 : _GEN_341;
  assign _GEN_343 = 10'h157 == index ? 32'h3000000 : _GEN_342;
  assign _GEN_344 = 10'h158 == index ? 32'h8000000 : _GEN_343;
  assign _GEN_345 = 10'h159 == index ? 32'h24010000 : _GEN_344;
  assign _GEN_346 = 10'h15a == index ? 32'h1000000 : _GEN_345;
  assign _GEN_347 = 10'h15b == index ? 32'h2000000 : _GEN_346;
  assign _GEN_348 = 10'h15c == index ? 32'h2000000 : _GEN_347;
  assign _GEN_349 = 10'h15d == index ? 32'h1000000 : _GEN_348;
  assign _GEN_350 = 10'h15e == index ? 32'h65746e69 : _GEN_349;
  assign _GEN_351 = 10'h15f == index ? 32'h70757272 : _GEN_350;
  assign _GEN_352 = 10'h160 == index ? 32'h6f632d74 : _GEN_351;
  assign _GEN_353 = 10'h161 == index ? 32'h6f72746e : _GEN_352;
  assign _GEN_354 = 10'h162 == index ? 32'h72656c6c : _GEN_353;
  assign _GEN_355 = 10'h163 == index ? 32'h30306340 : _GEN_354;
  assign _GEN_356 = 10'h164 == index ? 32'h30303030 : _GEN_355;
  assign _GEN_357 = 10'h165 == index ? 32'h0 : _GEN_356;
  assign _GEN_358 = 10'h166 == index ? 32'h3000000 : _GEN_357;
  assign _GEN_359 = 10'h167 == index ? 32'h4000000 : _GEN_358;
  assign _GEN_360 = 10'h168 == index ? 32'hba000000 : _GEN_359;
  assign _GEN_361 = 10'h169 == index ? 32'h1000000 : _GEN_360;
  assign _GEN_362 = 10'h16a == index ? 32'h3000000 : _GEN_361;
  assign _GEN_363 = 10'h16b == index ? 32'hc000000 : _GEN_362;
  assign _GEN_364 = 10'h16c == index ? 32'h1b000000 : _GEN_363;
  assign _GEN_365 = 10'h16d == index ? 32'h63736972 : _GEN_364;
  assign _GEN_366 = 10'h16e == index ? 32'h6c702c76 : _GEN_365;
  assign _GEN_367 = 10'h16f == index ? 32'h306369 : _GEN_366;
  assign _GEN_368 = 10'h170 == index ? 32'h3000000 : _GEN_367;
  assign _GEN_369 = 10'h171 == index ? 32'h0 : _GEN_368;
  assign _GEN_370 = 10'h172 == index ? 32'hcb000000 : _GEN_369;
  assign _GEN_371 = 10'h173 == index ? 32'h3000000 : _GEN_370;
  assign _GEN_372 = 10'h174 == index ? 32'h8000000 : _GEN_371;
  assign _GEN_373 = 10'h175 == index ? 32'hf5000000 : _GEN_372;
  assign _GEN_374 = 10'h176 == index ? 32'h3000000 : _GEN_373;
  assign _GEN_375 = 10'h177 == index ? 32'hb000000 : _GEN_374;
  assign _GEN_376 = 10'h178 == index ? 32'h3000000 : _GEN_375;
  assign _GEN_377 = 10'h179 == index ? 32'h8000000 : _GEN_376;
  assign _GEN_378 = 10'h17a == index ? 32'h99000000 : _GEN_377;
  assign _GEN_379 = 10'h17b == index ? 32'hc : _GEN_378;
  assign _GEN_380 = 10'h17c == index ? 32'h4 : _GEN_379;
  assign _GEN_381 = 10'h17d == index ? 32'h3000000 : _GEN_380;
  assign _GEN_382 = 10'h17e == index ? 32'h8000000 : _GEN_381;
  assign _GEN_383 = 10'h17f == index ? 32'h9010000 : _GEN_382;
  assign _GEN_384 = 10'h180 == index ? 32'h746e6f63 : _GEN_383;
  assign _GEN_385 = 10'h181 == index ? 32'h6c6f72 : _GEN_384;
  assign _GEN_386 = 10'h182 == index ? 32'h3000000 : _GEN_385;
  assign _GEN_387 = 10'h183 == index ? 32'h4000000 : _GEN_386;
  assign _GEN_388 = 10'h184 == index ? 32'h2f010000 : _GEN_387;
  assign _GEN_389 = 10'h185 == index ? 32'h7000000 : _GEN_388;
  assign _GEN_390 = 10'h186 == index ? 32'h3000000 : _GEN_389;
  assign _GEN_391 = 10'h187 == index ? 32'h4000000 : _GEN_390;
  assign _GEN_392 = 10'h188 == index ? 32'h42010000 : _GEN_391;
  assign _GEN_393 = 10'h189 == index ? 32'h2000000 : _GEN_392;
  assign _GEN_394 = 10'h18a == index ? 32'h3000000 : _GEN_393;
  assign _GEN_395 = 10'h18b == index ? 32'h4000000 : _GEN_394;
  assign _GEN_396 = 10'h18c == index ? 32'he0000000 : _GEN_395;
  assign _GEN_397 = 10'h18d == index ? 32'h4000000 : _GEN_396;
  assign _GEN_398 = 10'h18e == index ? 32'h3000000 : _GEN_397;
  assign _GEN_399 = 10'h18f == index ? 32'h4000000 : _GEN_398;
  assign _GEN_400 = 10'h190 == index ? 32'he6000000 : _GEN_399;
  assign _GEN_401 = 10'h191 == index ? 32'h4000000 : _GEN_400;
  assign _GEN_402 = 10'h192 == index ? 32'h2000000 : _GEN_401;
  assign _GEN_403 = 10'h193 == index ? 32'h1000000 : _GEN_402;
  assign _GEN_404 = 10'h194 == index ? 32'h6f696d6d : _GEN_403;
  assign _GEN_405 = 10'h195 == index ? 32'h30303640 : _GEN_404;
  assign _GEN_406 = 10'h196 == index ? 32'h30303030 : _GEN_405;
  assign _GEN_407 = 10'h197 == index ? 32'h30 : _GEN_406;
  assign _GEN_408 = 10'h198 == index ? 32'h3000000 : _GEN_407;
  assign _GEN_409 = 10'h199 == index ? 32'h4000000 : _GEN_408;
  assign _GEN_410 = 10'h19a == index ? 32'h0 : _GEN_409;
  assign _GEN_411 = 10'h19b == index ? 32'h1000000 : _GEN_410;
  assign _GEN_412 = 10'h19c == index ? 32'h3000000 : _GEN_411;
  assign _GEN_413 = 10'h19d == index ? 32'h4000000 : _GEN_412;
  assign _GEN_414 = 10'h19e == index ? 32'hf000000 : _GEN_413;
  assign _GEN_415 = 10'h19f == index ? 32'h1000000 : _GEN_414;
  assign _GEN_416 = 10'h1a0 == index ? 32'h3000000 : _GEN_415;
  assign _GEN_417 = 10'h1a1 == index ? 32'hb000000 : _GEN_416;
  assign _GEN_418 = 10'h1a2 == index ? 32'h1b000000 : _GEN_417;
  assign _GEN_419 = 10'h1a3 == index ? 32'h706d6973 : _GEN_418;
  assign _GEN_420 = 10'h1a4 == index ? 32'h622d656c : _GEN_419;
  assign _GEN_421 = 10'h1a5 == index ? 32'h7375 : _GEN_420;
  assign _GEN_422 = 10'h1a6 == index ? 32'h3000000 : _GEN_421;
  assign _GEN_423 = 10'h1a7 == index ? 32'hc000000 : _GEN_422;
  assign _GEN_424 = 10'h1a8 == index ? 32'hee000000 : _GEN_423;
  assign _GEN_425 = 10'h1a9 == index ? 32'h60 : _GEN_424;
  assign _GEN_426 = 10'h1aa == index ? 32'h60 : _GEN_425;
  assign _GEN_427 = 10'h1ab == index ? 32'h20 : _GEN_426;
  assign _GEN_428 = 10'h1ac == index ? 32'h2000000 : _GEN_427;
  assign _GEN_429 = 10'h1ad == index ? 32'h1000000 : _GEN_428;
  assign _GEN_430 = 10'h1ae == index ? 32'h406d6f72 : _GEN_429;
  assign _GEN_431 = 10'h1af == index ? 32'h30303031 : _GEN_430;
  assign _GEN_432 = 10'h1b0 == index ? 32'h30 : _GEN_431;
  assign _GEN_433 = 10'h1b1 == index ? 32'h3000000 : _GEN_432;
  assign _GEN_434 = 10'h1b2 == index ? 32'hc000000 : _GEN_433;
  assign _GEN_435 = 10'h1b3 == index ? 32'h1b000000 : _GEN_434;
  assign _GEN_436 = 10'h1b4 == index ? 32'h69666973 : _GEN_435;
  assign _GEN_437 = 10'h1b5 == index ? 32'h722c6576 : _GEN_436;
  assign _GEN_438 = 10'h1b6 == index ? 32'h306d6f : _GEN_437;
  assign _GEN_439 = 10'h1b7 == index ? 32'h3000000 : _GEN_438;
  assign _GEN_440 = 10'h1b8 == index ? 32'h8000000 : _GEN_439;
  assign _GEN_441 = 10'h1b9 == index ? 32'h99000000 : _GEN_440;
  assign _GEN_442 = 10'h1ba == index ? 32'h100 : _GEN_441;
  assign _GEN_443 = 10'h1bb == index ? 32'h100 : _GEN_442;
  assign _GEN_444 = 10'h1bc == index ? 32'h3000000 : _GEN_443;
  assign _GEN_445 = 10'h1bd == index ? 32'h4000000 : _GEN_444;
  assign _GEN_446 = 10'h1be == index ? 32'h9010000 : _GEN_445;
  assign _GEN_447 = 10'h1bf == index ? 32'h6d656d : _GEN_446;
  assign _GEN_448 = 10'h1c0 == index ? 32'h2000000 : _GEN_447;
  assign _GEN_449 = 10'h1c1 == index ? 32'h2000000 : _GEN_448;
  assign _GEN_450 = 10'h1c2 == index ? 32'h2000000 : _GEN_449;
  assign _GEN_451 = 10'h1c3 == index ? 32'h9000000 : _GEN_450;
  assign _GEN_452 = 10'h1c4 == index ? 32'h64646123 : _GEN_451;
  assign _GEN_453 = 10'h1c5 == index ? 32'h73736572 : _GEN_452;
  assign _GEN_454 = 10'h1c6 == index ? 32'h6c65632d : _GEN_453;
  assign _GEN_455 = 10'h1c7 == index ? 32'h2300736c : _GEN_454;
  assign _GEN_456 = 10'h1c8 == index ? 32'h657a6973 : _GEN_455;
  assign _GEN_457 = 10'h1c9 == index ? 32'h6c65632d : _GEN_456;
  assign _GEN_458 = 10'h1ca == index ? 32'h6300736c : _GEN_457;
  assign _GEN_459 = 10'h1cb == index ? 32'h61706d6f : _GEN_458;
  assign _GEN_460 = 10'h1cc == index ? 32'h6c626974 : _GEN_459;
  assign _GEN_461 = 10'h1cd == index ? 32'h6f6d0065 : _GEN_460;
  assign _GEN_462 = 10'h1ce == index ? 32'h6c6564 : _GEN_461;
  assign _GEN_463 = 10'h1cf == index ? 32'h656d6974 : _GEN_462;
  assign _GEN_464 = 10'h1d0 == index ? 32'h65736162 : _GEN_463;
  assign _GEN_465 = 10'h1d1 == index ? 32'h6572662d : _GEN_464;
  assign _GEN_466 = 10'h1d2 == index ? 32'h6e657571 : _GEN_465;
  assign _GEN_467 = 10'h1d3 == index ? 32'h63007963 : _GEN_466;
  assign _GEN_468 = 10'h1d4 == index ? 32'h6b636f6c : _GEN_467;
  assign _GEN_469 = 10'h1d5 == index ? 32'h6572662d : _GEN_468;
  assign _GEN_470 = 10'h1d6 == index ? 32'h6e657571 : _GEN_469;
  assign _GEN_471 = 10'h1d7 == index ? 32'h64007963 : _GEN_470;
  assign _GEN_472 = 10'h1d8 == index ? 32'h63697665 : _GEN_471;
  assign _GEN_473 = 10'h1d9 == index ? 32'h79745f65 : _GEN_472;
  assign _GEN_474 = 10'h1da == index ? 32'h69006570 : _GEN_473;
  assign _GEN_475 = 10'h1db == index ? 32'h6361632d : _GEN_474;
  assign _GEN_476 = 10'h1dc == index ? 32'h622d6568 : _GEN_475;
  assign _GEN_477 = 10'h1dd == index ? 32'h6b636f6c : _GEN_476;
  assign _GEN_478 = 10'h1de == index ? 32'h7a69732d : _GEN_477;
  assign _GEN_479 = 10'h1df == index ? 32'h2d690065 : _GEN_478;
  assign _GEN_480 = 10'h1e0 == index ? 32'h68636163 : _GEN_479;
  assign _GEN_481 = 10'h1e1 == index ? 32'h65732d65 : _GEN_480;
  assign _GEN_482 = 10'h1e2 == index ? 32'h69007374 : _GEN_481;
  assign _GEN_483 = 10'h1e3 == index ? 32'h6361632d : _GEN_482;
  assign _GEN_484 = 10'h1e4 == index ? 32'h732d6568 : _GEN_483;
  assign _GEN_485 = 10'h1e5 == index ? 32'h657a69 : _GEN_484;
  assign _GEN_486 = 10'h1e6 == index ? 32'h7478656e : _GEN_485;
  assign _GEN_487 = 10'h1e7 == index ? 32'h76656c2d : _GEN_486;
  assign _GEN_488 = 10'h1e8 == index ? 32'h632d6c65 : _GEN_487;
  assign _GEN_489 = 10'h1e9 == index ? 32'h65686361 : _GEN_488;
  assign _GEN_490 = 10'h1ea == index ? 32'h67657200 : _GEN_489;
  assign _GEN_491 = 10'h1eb == index ? 32'h73697200 : _GEN_490;
  assign _GEN_492 = 10'h1ec == index ? 32'h692c7663 : _GEN_491;
  assign _GEN_493 = 10'h1ed == index ? 32'h73006173 : _GEN_492;
  assign _GEN_494 = 10'h1ee == index ? 32'h76696669 : _GEN_493;
  assign _GEN_495 = 10'h1ef == index ? 32'h74642c65 : _GEN_494;
  assign _GEN_496 = 10'h1f0 == index ? 32'h73006d69 : _GEN_495;
  assign _GEN_497 = 10'h1f1 == index ? 32'h75746174 : _GEN_496;
  assign _GEN_498 = 10'h1f2 == index ? 32'h69230073 : _GEN_497;
  assign _GEN_499 = 10'h1f3 == index ? 32'h7265746e : _GEN_498;
  assign _GEN_500 = 10'h1f4 == index ? 32'h74707572 : _GEN_499;
  assign _GEN_501 = 10'h1f5 == index ? 32'h6c65632d : _GEN_500;
  assign _GEN_502 = 10'h1f6 == index ? 32'h6900736c : _GEN_501;
  assign _GEN_503 = 10'h1f7 == index ? 32'h7265746e : _GEN_502;
  assign _GEN_504 = 10'h1f8 == index ? 32'h74707572 : _GEN_503;
  assign _GEN_505 = 10'h1f9 == index ? 32'h6e6f632d : _GEN_504;
  assign _GEN_506 = 10'h1fa == index ? 32'h6c6f7274 : _GEN_505;
  assign _GEN_507 = 10'h1fb == index ? 32'h72656c : _GEN_506;
  assign _GEN_508 = 10'h1fc == index ? 32'h756e696c : _GEN_507;
  assign _GEN_509 = 10'h1fd == index ? 32'h68702c78 : _GEN_508;
  assign _GEN_510 = 10'h1fe == index ? 32'h6c646e61 : _GEN_509;
  assign _GEN_511 = 10'h1ff == index ? 32'h61720065 : _GEN_510;
  assign _GEN_512 = 10'h200 == index ? 32'h7365676e : _GEN_511;
  assign _GEN_513 = 10'h201 == index ? 32'h746e6900 : _GEN_512;
  assign _GEN_514 = 10'h202 == index ? 32'h75727265 : _GEN_513;
  assign _GEN_515 = 10'h203 == index ? 32'h2d737470 : _GEN_514;
  assign _GEN_516 = 10'h204 == index ? 32'h65747865 : _GEN_515;
  assign _GEN_517 = 10'h205 == index ? 32'h6465646e : _GEN_516;
  assign _GEN_518 = 10'h206 == index ? 32'h67657200 : _GEN_517;
  assign _GEN_519 = 10'h207 == index ? 32'h6d616e2d : _GEN_518;
  assign _GEN_520 = 10'h208 == index ? 32'h69007365 : _GEN_519;
  assign _GEN_521 = 10'h209 == index ? 32'h7265746e : _GEN_520;
  assign _GEN_522 = 10'h20a == index ? 32'h74707572 : _GEN_521;
  assign _GEN_523 = 10'h20b == index ? 32'h7261702d : _GEN_522;
  assign _GEN_524 = 10'h20c == index ? 32'h746e65 : _GEN_523;
  assign _GEN_525 = 10'h20d == index ? 32'h65746e69 : _GEN_524;
  assign _GEN_526 = 10'h20e == index ? 32'h70757272 : _GEN_525;
  assign _GEN_527 = 10'h20f == index ? 32'h72007374 : _GEN_526;
  assign _GEN_528 = 10'h210 == index ? 32'h76637369 : _GEN_527;
  assign _GEN_529 = 10'h211 == index ? 32'h78616d2c : _GEN_528;
  assign _GEN_530 = 10'h212 == index ? 32'h6972702d : _GEN_529;
  assign _GEN_531 = 10'h213 == index ? 32'h7469726f : _GEN_530;
  assign _GEN_532 = 10'h214 == index ? 32'h69720079 : _GEN_531;
  assign _GEN_533 = 10'h215 == index ? 32'h2c766373 : _GEN_532;
  assign _GEN_534 = 10'h216 == index ? 32'h7665646e : _GEN_533;
  assign _GEN_535 = 10'h217 == index ? 32'h0 : _GEN_534;
  assign _GEN_536 = 10'h218 == index ? 32'h0 : _GEN_535;
  assign _GEN_537 = 10'h219 == index ? 32'h0 : _GEN_536;
  assign _GEN_538 = 10'h21a == index ? 32'h0 : _GEN_537;
  assign _GEN_539 = 10'h21b == index ? 32'h0 : _GEN_538;
  assign _GEN_540 = 10'h21c == index ? 32'h0 : _GEN_539;
  assign _GEN_541 = 10'h21d == index ? 32'h0 : _GEN_540;
  assign _GEN_542 = 10'h21e == index ? 32'h0 : _GEN_541;
  assign _GEN_543 = 10'h21f == index ? 32'h0 : _GEN_542;
  assign _GEN_544 = 10'h220 == index ? 32'h0 : _GEN_543;
  assign _GEN_545 = 10'h221 == index ? 32'h0 : _GEN_544;
  assign _GEN_546 = 10'h222 == index ? 32'h0 : _GEN_545;
  assign _GEN_547 = 10'h223 == index ? 32'h0 : _GEN_546;
  assign _GEN_548 = 10'h224 == index ? 32'h0 : _GEN_547;
  assign _GEN_549 = 10'h225 == index ? 32'h0 : _GEN_548;
  assign _GEN_550 = 10'h226 == index ? 32'h0 : _GEN_549;
  assign _GEN_551 = 10'h227 == index ? 32'h0 : _GEN_550;
  assign _GEN_552 = 10'h228 == index ? 32'h0 : _GEN_551;
  assign _GEN_553 = 10'h229 == index ? 32'h0 : _GEN_552;
  assign _GEN_554 = 10'h22a == index ? 32'h0 : _GEN_553;
  assign _GEN_555 = 10'h22b == index ? 32'h0 : _GEN_554;
  assign _GEN_556 = 10'h22c == index ? 32'h0 : _GEN_555;
  assign _GEN_557 = 10'h22d == index ? 32'h0 : _GEN_556;
  assign _GEN_558 = 10'h22e == index ? 32'h0 : _GEN_557;
  assign _GEN_559 = 10'h22f == index ? 32'h0 : _GEN_558;
  assign _GEN_560 = 10'h230 == index ? 32'h0 : _GEN_559;
  assign _GEN_561 = 10'h231 == index ? 32'h0 : _GEN_560;
  assign _GEN_562 = 10'h232 == index ? 32'h0 : _GEN_561;
  assign _GEN_563 = 10'h233 == index ? 32'h0 : _GEN_562;
  assign _GEN_564 = 10'h234 == index ? 32'h0 : _GEN_563;
  assign _GEN_565 = 10'h235 == index ? 32'h0 : _GEN_564;
  assign _GEN_566 = 10'h236 == index ? 32'h0 : _GEN_565;
  assign _GEN_567 = 10'h237 == index ? 32'h0 : _GEN_566;
  assign _GEN_568 = 10'h238 == index ? 32'h0 : _GEN_567;
  assign _GEN_569 = 10'h239 == index ? 32'h0 : _GEN_568;
  assign _GEN_570 = 10'h23a == index ? 32'h0 : _GEN_569;
  assign _GEN_571 = 10'h23b == index ? 32'h0 : _GEN_570;
  assign _GEN_572 = 10'h23c == index ? 32'h0 : _GEN_571;
  assign _GEN_573 = 10'h23d == index ? 32'h0 : _GEN_572;
  assign _GEN_574 = 10'h23e == index ? 32'h0 : _GEN_573;
  assign _GEN_575 = 10'h23f == index ? 32'h0 : _GEN_574;
  assign _GEN_576 = 10'h240 == index ? 32'h0 : _GEN_575;
  assign _GEN_577 = 10'h241 == index ? 32'h0 : _GEN_576;
  assign _GEN_578 = 10'h242 == index ? 32'h0 : _GEN_577;
  assign _GEN_579 = 10'h243 == index ? 32'h0 : _GEN_578;
  assign _GEN_580 = 10'h244 == index ? 32'h0 : _GEN_579;
  assign _GEN_581 = 10'h245 == index ? 32'h0 : _GEN_580;
  assign _GEN_582 = 10'h246 == index ? 32'h0 : _GEN_581;
  assign _GEN_583 = 10'h247 == index ? 32'h0 : _GEN_582;
  assign _GEN_584 = 10'h248 == index ? 32'h0 : _GEN_583;
  assign _GEN_585 = 10'h249 == index ? 32'h0 : _GEN_584;
  assign _GEN_586 = 10'h24a == index ? 32'h0 : _GEN_585;
  assign _GEN_587 = 10'h24b == index ? 32'h0 : _GEN_586;
  assign _GEN_588 = 10'h24c == index ? 32'h0 : _GEN_587;
  assign _GEN_589 = 10'h24d == index ? 32'h0 : _GEN_588;
  assign _GEN_590 = 10'h24e == index ? 32'h0 : _GEN_589;
  assign _GEN_591 = 10'h24f == index ? 32'h0 : _GEN_590;
  assign _GEN_592 = 10'h250 == index ? 32'h0 : _GEN_591;
  assign _GEN_593 = 10'h251 == index ? 32'h0 : _GEN_592;
  assign _GEN_594 = 10'h252 == index ? 32'h0 : _GEN_593;
  assign _GEN_595 = 10'h253 == index ? 32'h0 : _GEN_594;
  assign _GEN_596 = 10'h254 == index ? 32'h0 : _GEN_595;
  assign _GEN_597 = 10'h255 == index ? 32'h0 : _GEN_596;
  assign _GEN_598 = 10'h256 == index ? 32'h0 : _GEN_597;
  assign _GEN_599 = 10'h257 == index ? 32'h0 : _GEN_598;
  assign _GEN_600 = 10'h258 == index ? 32'h0 : _GEN_599;
  assign _GEN_601 = 10'h259 == index ? 32'h0 : _GEN_600;
  assign _GEN_602 = 10'h25a == index ? 32'h0 : _GEN_601;
  assign _GEN_603 = 10'h25b == index ? 32'h0 : _GEN_602;
  assign _GEN_604 = 10'h25c == index ? 32'h0 : _GEN_603;
  assign _GEN_605 = 10'h25d == index ? 32'h0 : _GEN_604;
  assign _GEN_606 = 10'h25e == index ? 32'h0 : _GEN_605;
  assign _GEN_607 = 10'h25f == index ? 32'h0 : _GEN_606;
  assign _GEN_608 = 10'h260 == index ? 32'h0 : _GEN_607;
  assign _GEN_609 = 10'h261 == index ? 32'h0 : _GEN_608;
  assign _GEN_610 = 10'h262 == index ? 32'h0 : _GEN_609;
  assign _GEN_611 = 10'h263 == index ? 32'h0 : _GEN_610;
  assign _GEN_612 = 10'h264 == index ? 32'h0 : _GEN_611;
  assign _GEN_613 = 10'h265 == index ? 32'h0 : _GEN_612;
  assign _GEN_614 = 10'h266 == index ? 32'h0 : _GEN_613;
  assign _GEN_615 = 10'h267 == index ? 32'h0 : _GEN_614;
  assign _GEN_616 = 10'h268 == index ? 32'h0 : _GEN_615;
  assign _GEN_617 = 10'h269 == index ? 32'h0 : _GEN_616;
  assign _GEN_618 = 10'h26a == index ? 32'h0 : _GEN_617;
  assign _GEN_619 = 10'h26b == index ? 32'h0 : _GEN_618;
  assign _GEN_620 = 10'h26c == index ? 32'h0 : _GEN_619;
  assign _GEN_621 = 10'h26d == index ? 32'h0 : _GEN_620;
  assign _GEN_622 = 10'h26e == index ? 32'h0 : _GEN_621;
  assign _GEN_623 = 10'h26f == index ? 32'h0 : _GEN_622;
  assign _GEN_624 = 10'h270 == index ? 32'h0 : _GEN_623;
  assign _GEN_625 = 10'h271 == index ? 32'h0 : _GEN_624;
  assign _GEN_626 = 10'h272 == index ? 32'h0 : _GEN_625;
  assign _GEN_627 = 10'h273 == index ? 32'h0 : _GEN_626;
  assign _GEN_628 = 10'h274 == index ? 32'h0 : _GEN_627;
  assign _GEN_629 = 10'h275 == index ? 32'h0 : _GEN_628;
  assign _GEN_630 = 10'h276 == index ? 32'h0 : _GEN_629;
  assign _GEN_631 = 10'h277 == index ? 32'h0 : _GEN_630;
  assign _GEN_632 = 10'h278 == index ? 32'h0 : _GEN_631;
  assign _GEN_633 = 10'h279 == index ? 32'h0 : _GEN_632;
  assign _GEN_634 = 10'h27a == index ? 32'h0 : _GEN_633;
  assign _GEN_635 = 10'h27b == index ? 32'h0 : _GEN_634;
  assign _GEN_636 = 10'h27c == index ? 32'h0 : _GEN_635;
  assign _GEN_637 = 10'h27d == index ? 32'h0 : _GEN_636;
  assign _GEN_638 = 10'h27e == index ? 32'h0 : _GEN_637;
  assign _GEN_639 = 10'h27f == index ? 32'h0 : _GEN_638;
  assign _GEN_640 = 10'h280 == index ? 32'h0 : _GEN_639;
  assign _GEN_641 = 10'h281 == index ? 32'h0 : _GEN_640;
  assign _GEN_642 = 10'h282 == index ? 32'h0 : _GEN_641;
  assign _GEN_643 = 10'h283 == index ? 32'h0 : _GEN_642;
  assign _GEN_644 = 10'h284 == index ? 32'h0 : _GEN_643;
  assign _GEN_645 = 10'h285 == index ? 32'h0 : _GEN_644;
  assign _GEN_646 = 10'h286 == index ? 32'h0 : _GEN_645;
  assign _GEN_647 = 10'h287 == index ? 32'h0 : _GEN_646;
  assign _GEN_648 = 10'h288 == index ? 32'h0 : _GEN_647;
  assign _GEN_649 = 10'h289 == index ? 32'h0 : _GEN_648;
  assign _GEN_650 = 10'h28a == index ? 32'h0 : _GEN_649;
  assign _GEN_651 = 10'h28b == index ? 32'h0 : _GEN_650;
  assign _GEN_652 = 10'h28c == index ? 32'h0 : _GEN_651;
  assign _GEN_653 = 10'h28d == index ? 32'h0 : _GEN_652;
  assign _GEN_654 = 10'h28e == index ? 32'h0 : _GEN_653;
  assign _GEN_655 = 10'h28f == index ? 32'h0 : _GEN_654;
  assign _GEN_656 = 10'h290 == index ? 32'h0 : _GEN_655;
  assign _GEN_657 = 10'h291 == index ? 32'h0 : _GEN_656;
  assign _GEN_658 = 10'h292 == index ? 32'h0 : _GEN_657;
  assign _GEN_659 = 10'h293 == index ? 32'h0 : _GEN_658;
  assign _GEN_660 = 10'h294 == index ? 32'h0 : _GEN_659;
  assign _GEN_661 = 10'h295 == index ? 32'h0 : _GEN_660;
  assign _GEN_662 = 10'h296 == index ? 32'h0 : _GEN_661;
  assign _GEN_663 = 10'h297 == index ? 32'h0 : _GEN_662;
  assign _GEN_664 = 10'h298 == index ? 32'h0 : _GEN_663;
  assign _GEN_665 = 10'h299 == index ? 32'h0 : _GEN_664;
  assign _GEN_666 = 10'h29a == index ? 32'h0 : _GEN_665;
  assign _GEN_667 = 10'h29b == index ? 32'h0 : _GEN_666;
  assign _GEN_668 = 10'h29c == index ? 32'h0 : _GEN_667;
  assign _GEN_669 = 10'h29d == index ? 32'h0 : _GEN_668;
  assign _GEN_670 = 10'h29e == index ? 32'h0 : _GEN_669;
  assign _GEN_671 = 10'h29f == index ? 32'h0 : _GEN_670;
  assign _GEN_672 = 10'h2a0 == index ? 32'h0 : _GEN_671;
  assign _GEN_673 = 10'h2a1 == index ? 32'h0 : _GEN_672;
  assign _GEN_674 = 10'h2a2 == index ? 32'h0 : _GEN_673;
  assign _GEN_675 = 10'h2a3 == index ? 32'h0 : _GEN_674;
  assign _GEN_676 = 10'h2a4 == index ? 32'h0 : _GEN_675;
  assign _GEN_677 = 10'h2a5 == index ? 32'h0 : _GEN_676;
  assign _GEN_678 = 10'h2a6 == index ? 32'h0 : _GEN_677;
  assign _GEN_679 = 10'h2a7 == index ? 32'h0 : _GEN_678;
  assign _GEN_680 = 10'h2a8 == index ? 32'h0 : _GEN_679;
  assign _GEN_681 = 10'h2a9 == index ? 32'h0 : _GEN_680;
  assign _GEN_682 = 10'h2aa == index ? 32'h0 : _GEN_681;
  assign _GEN_683 = 10'h2ab == index ? 32'h0 : _GEN_682;
  assign _GEN_684 = 10'h2ac == index ? 32'h0 : _GEN_683;
  assign _GEN_685 = 10'h2ad == index ? 32'h0 : _GEN_684;
  assign _GEN_686 = 10'h2ae == index ? 32'h0 : _GEN_685;
  assign _GEN_687 = 10'h2af == index ? 32'h0 : _GEN_686;
  assign _GEN_688 = 10'h2b0 == index ? 32'h0 : _GEN_687;
  assign _GEN_689 = 10'h2b1 == index ? 32'h0 : _GEN_688;
  assign _GEN_690 = 10'h2b2 == index ? 32'h0 : _GEN_689;
  assign _GEN_691 = 10'h2b3 == index ? 32'h0 : _GEN_690;
  assign _GEN_692 = 10'h2b4 == index ? 32'h0 : _GEN_691;
  assign _GEN_693 = 10'h2b5 == index ? 32'h0 : _GEN_692;
  assign _GEN_694 = 10'h2b6 == index ? 32'h0 : _GEN_693;
  assign _GEN_695 = 10'h2b7 == index ? 32'h0 : _GEN_694;
  assign _GEN_696 = 10'h2b8 == index ? 32'h0 : _GEN_695;
  assign _GEN_697 = 10'h2b9 == index ? 32'h0 : _GEN_696;
  assign _GEN_698 = 10'h2ba == index ? 32'h0 : _GEN_697;
  assign _GEN_699 = 10'h2bb == index ? 32'h0 : _GEN_698;
  assign _GEN_700 = 10'h2bc == index ? 32'h0 : _GEN_699;
  assign _GEN_701 = 10'h2bd == index ? 32'h0 : _GEN_700;
  assign _GEN_702 = 10'h2be == index ? 32'h0 : _GEN_701;
  assign _GEN_703 = 10'h2bf == index ? 32'h0 : _GEN_702;
  assign _GEN_704 = 10'h2c0 == index ? 32'h0 : _GEN_703;
  assign _GEN_705 = 10'h2c1 == index ? 32'h0 : _GEN_704;
  assign _GEN_706 = 10'h2c2 == index ? 32'h0 : _GEN_705;
  assign _GEN_707 = 10'h2c3 == index ? 32'h0 : _GEN_706;
  assign _GEN_708 = 10'h2c4 == index ? 32'h0 : _GEN_707;
  assign _GEN_709 = 10'h2c5 == index ? 32'h0 : _GEN_708;
  assign _GEN_710 = 10'h2c6 == index ? 32'h0 : _GEN_709;
  assign _GEN_711 = 10'h2c7 == index ? 32'h0 : _GEN_710;
  assign _GEN_712 = 10'h2c8 == index ? 32'h0 : _GEN_711;
  assign _GEN_713 = 10'h2c9 == index ? 32'h0 : _GEN_712;
  assign _GEN_714 = 10'h2ca == index ? 32'h0 : _GEN_713;
  assign _GEN_715 = 10'h2cb == index ? 32'h0 : _GEN_714;
  assign _GEN_716 = 10'h2cc == index ? 32'h0 : _GEN_715;
  assign _GEN_717 = 10'h2cd == index ? 32'h0 : _GEN_716;
  assign _GEN_718 = 10'h2ce == index ? 32'h0 : _GEN_717;
  assign _GEN_719 = 10'h2cf == index ? 32'h0 : _GEN_718;
  assign _GEN_720 = 10'h2d0 == index ? 32'h0 : _GEN_719;
  assign _GEN_721 = 10'h2d1 == index ? 32'h0 : _GEN_720;
  assign _GEN_722 = 10'h2d2 == index ? 32'h0 : _GEN_721;
  assign _GEN_723 = 10'h2d3 == index ? 32'h0 : _GEN_722;
  assign _GEN_724 = 10'h2d4 == index ? 32'h0 : _GEN_723;
  assign _GEN_725 = 10'h2d5 == index ? 32'h0 : _GEN_724;
  assign _GEN_726 = 10'h2d6 == index ? 32'h0 : _GEN_725;
  assign _GEN_727 = 10'h2d7 == index ? 32'h0 : _GEN_726;
  assign _GEN_728 = 10'h2d8 == index ? 32'h0 : _GEN_727;
  assign _GEN_729 = 10'h2d9 == index ? 32'h0 : _GEN_728;
  assign _GEN_730 = 10'h2da == index ? 32'h0 : _GEN_729;
  assign _GEN_731 = 10'h2db == index ? 32'h0 : _GEN_730;
  assign _GEN_732 = 10'h2dc == index ? 32'h0 : _GEN_731;
  assign _GEN_733 = 10'h2dd == index ? 32'h0 : _GEN_732;
  assign _GEN_734 = 10'h2de == index ? 32'h0 : _GEN_733;
  assign _GEN_735 = 10'h2df == index ? 32'h0 : _GEN_734;
  assign _GEN_736 = 10'h2e0 == index ? 32'h0 : _GEN_735;
  assign _GEN_737 = 10'h2e1 == index ? 32'h0 : _GEN_736;
  assign _GEN_738 = 10'h2e2 == index ? 32'h0 : _GEN_737;
  assign _GEN_739 = 10'h2e3 == index ? 32'h0 : _GEN_738;
  assign _GEN_740 = 10'h2e4 == index ? 32'h0 : _GEN_739;
  assign _GEN_741 = 10'h2e5 == index ? 32'h0 : _GEN_740;
  assign _GEN_742 = 10'h2e6 == index ? 32'h0 : _GEN_741;
  assign _GEN_743 = 10'h2e7 == index ? 32'h0 : _GEN_742;
  assign _GEN_744 = 10'h2e8 == index ? 32'h0 : _GEN_743;
  assign _GEN_745 = 10'h2e9 == index ? 32'h0 : _GEN_744;
  assign _GEN_746 = 10'h2ea == index ? 32'h0 : _GEN_745;
  assign _GEN_747 = 10'h2eb == index ? 32'h0 : _GEN_746;
  assign _GEN_748 = 10'h2ec == index ? 32'h0 : _GEN_747;
  assign _GEN_749 = 10'h2ed == index ? 32'h0 : _GEN_748;
  assign _GEN_750 = 10'h2ee == index ? 32'h0 : _GEN_749;
  assign _GEN_751 = 10'h2ef == index ? 32'h0 : _GEN_750;
  assign _GEN_752 = 10'h2f0 == index ? 32'h0 : _GEN_751;
  assign _GEN_753 = 10'h2f1 == index ? 32'h0 : _GEN_752;
  assign _GEN_754 = 10'h2f2 == index ? 32'h0 : _GEN_753;
  assign _GEN_755 = 10'h2f3 == index ? 32'h0 : _GEN_754;
  assign _GEN_756 = 10'h2f4 == index ? 32'h0 : _GEN_755;
  assign _GEN_757 = 10'h2f5 == index ? 32'h0 : _GEN_756;
  assign _GEN_758 = 10'h2f6 == index ? 32'h0 : _GEN_757;
  assign _GEN_759 = 10'h2f7 == index ? 32'h0 : _GEN_758;
  assign _GEN_760 = 10'h2f8 == index ? 32'h0 : _GEN_759;
  assign _GEN_761 = 10'h2f9 == index ? 32'h0 : _GEN_760;
  assign _GEN_762 = 10'h2fa == index ? 32'h0 : _GEN_761;
  assign _GEN_763 = 10'h2fb == index ? 32'h0 : _GEN_762;
  assign _GEN_764 = 10'h2fc == index ? 32'h0 : _GEN_763;
  assign _GEN_765 = 10'h2fd == index ? 32'h0 : _GEN_764;
  assign _GEN_766 = 10'h2fe == index ? 32'h0 : _GEN_765;
  assign _GEN_767 = 10'h2ff == index ? 32'h0 : _GEN_766;
  assign _GEN_768 = 10'h300 == index ? 32'h0 : _GEN_767;
  assign _GEN_769 = 10'h301 == index ? 32'h0 : _GEN_768;
  assign _GEN_770 = 10'h302 == index ? 32'h0 : _GEN_769;
  assign _GEN_771 = 10'h303 == index ? 32'h0 : _GEN_770;
  assign _GEN_772 = 10'h304 == index ? 32'h0 : _GEN_771;
  assign _GEN_773 = 10'h305 == index ? 32'h0 : _GEN_772;
  assign _GEN_774 = 10'h306 == index ? 32'h0 : _GEN_773;
  assign _GEN_775 = 10'h307 == index ? 32'h0 : _GEN_774;
  assign _GEN_776 = 10'h308 == index ? 32'h0 : _GEN_775;
  assign _GEN_777 = 10'h309 == index ? 32'h0 : _GEN_776;
  assign _GEN_778 = 10'h30a == index ? 32'h0 : _GEN_777;
  assign _GEN_779 = 10'h30b == index ? 32'h0 : _GEN_778;
  assign _GEN_780 = 10'h30c == index ? 32'h0 : _GEN_779;
  assign _GEN_781 = 10'h30d == index ? 32'h0 : _GEN_780;
  assign _GEN_782 = 10'h30e == index ? 32'h0 : _GEN_781;
  assign _GEN_783 = 10'h30f == index ? 32'h0 : _GEN_782;
  assign _GEN_784 = 10'h310 == index ? 32'h0 : _GEN_783;
  assign _GEN_785 = 10'h311 == index ? 32'h0 : _GEN_784;
  assign _GEN_786 = 10'h312 == index ? 32'h0 : _GEN_785;
  assign _GEN_787 = 10'h313 == index ? 32'h0 : _GEN_786;
  assign _GEN_788 = 10'h314 == index ? 32'h0 : _GEN_787;
  assign _GEN_789 = 10'h315 == index ? 32'h0 : _GEN_788;
  assign _GEN_790 = 10'h316 == index ? 32'h0 : _GEN_789;
  assign _GEN_791 = 10'h317 == index ? 32'h0 : _GEN_790;
  assign _GEN_792 = 10'h318 == index ? 32'h0 : _GEN_791;
  assign _GEN_793 = 10'h319 == index ? 32'h0 : _GEN_792;
  assign _GEN_794 = 10'h31a == index ? 32'h0 : _GEN_793;
  assign _GEN_795 = 10'h31b == index ? 32'h0 : _GEN_794;
  assign _GEN_796 = 10'h31c == index ? 32'h0 : _GEN_795;
  assign _GEN_797 = 10'h31d == index ? 32'h0 : _GEN_796;
  assign _GEN_798 = 10'h31e == index ? 32'h0 : _GEN_797;
  assign _GEN_799 = 10'h31f == index ? 32'h0 : _GEN_798;
  assign _GEN_800 = 10'h320 == index ? 32'h0 : _GEN_799;
  assign _GEN_801 = 10'h321 == index ? 32'h0 : _GEN_800;
  assign _GEN_802 = 10'h322 == index ? 32'h0 : _GEN_801;
  assign _GEN_803 = 10'h323 == index ? 32'h0 : _GEN_802;
  assign _GEN_804 = 10'h324 == index ? 32'h0 : _GEN_803;
  assign _GEN_805 = 10'h325 == index ? 32'h0 : _GEN_804;
  assign _GEN_806 = 10'h326 == index ? 32'h0 : _GEN_805;
  assign _GEN_807 = 10'h327 == index ? 32'h0 : _GEN_806;
  assign _GEN_808 = 10'h328 == index ? 32'h0 : _GEN_807;
  assign _GEN_809 = 10'h329 == index ? 32'h0 : _GEN_808;
  assign _GEN_810 = 10'h32a == index ? 32'h0 : _GEN_809;
  assign _GEN_811 = 10'h32b == index ? 32'h0 : _GEN_810;
  assign _GEN_812 = 10'h32c == index ? 32'h0 : _GEN_811;
  assign _GEN_813 = 10'h32d == index ? 32'h0 : _GEN_812;
  assign _GEN_814 = 10'h32e == index ? 32'h0 : _GEN_813;
  assign _GEN_815 = 10'h32f == index ? 32'h0 : _GEN_814;
  assign _GEN_816 = 10'h330 == index ? 32'h0 : _GEN_815;
  assign _GEN_817 = 10'h331 == index ? 32'h0 : _GEN_816;
  assign _GEN_818 = 10'h332 == index ? 32'h0 : _GEN_817;
  assign _GEN_819 = 10'h333 == index ? 32'h0 : _GEN_818;
  assign _GEN_820 = 10'h334 == index ? 32'h0 : _GEN_819;
  assign _GEN_821 = 10'h335 == index ? 32'h0 : _GEN_820;
  assign _GEN_822 = 10'h336 == index ? 32'h0 : _GEN_821;
  assign _GEN_823 = 10'h337 == index ? 32'h0 : _GEN_822;
  assign _GEN_824 = 10'h338 == index ? 32'h0 : _GEN_823;
  assign _GEN_825 = 10'h339 == index ? 32'h0 : _GEN_824;
  assign _GEN_826 = 10'h33a == index ? 32'h0 : _GEN_825;
  assign _GEN_827 = 10'h33b == index ? 32'h0 : _GEN_826;
  assign _GEN_828 = 10'h33c == index ? 32'h0 : _GEN_827;
  assign _GEN_829 = 10'h33d == index ? 32'h0 : _GEN_828;
  assign _GEN_830 = 10'h33e == index ? 32'h0 : _GEN_829;
  assign _GEN_831 = 10'h33f == index ? 32'h0 : _GEN_830;
  assign _GEN_832 = 10'h340 == index ? 32'h0 : _GEN_831;
  assign _GEN_833 = 10'h341 == index ? 32'h0 : _GEN_832;
  assign _GEN_834 = 10'h342 == index ? 32'h0 : _GEN_833;
  assign _GEN_835 = 10'h343 == index ? 32'h0 : _GEN_834;
  assign _GEN_836 = 10'h344 == index ? 32'h0 : _GEN_835;
  assign _GEN_837 = 10'h345 == index ? 32'h0 : _GEN_836;
  assign _GEN_838 = 10'h346 == index ? 32'h0 : _GEN_837;
  assign _GEN_839 = 10'h347 == index ? 32'h0 : _GEN_838;
  assign _GEN_840 = 10'h348 == index ? 32'h0 : _GEN_839;
  assign _GEN_841 = 10'h349 == index ? 32'h0 : _GEN_840;
  assign _GEN_842 = 10'h34a == index ? 32'h0 : _GEN_841;
  assign _GEN_843 = 10'h34b == index ? 32'h0 : _GEN_842;
  assign _GEN_844 = 10'h34c == index ? 32'h0 : _GEN_843;
  assign _GEN_845 = 10'h34d == index ? 32'h0 : _GEN_844;
  assign _GEN_846 = 10'h34e == index ? 32'h0 : _GEN_845;
  assign _GEN_847 = 10'h34f == index ? 32'h0 : _GEN_846;
  assign _GEN_848 = 10'h350 == index ? 32'h0 : _GEN_847;
  assign _GEN_849 = 10'h351 == index ? 32'h0 : _GEN_848;
  assign _GEN_850 = 10'h352 == index ? 32'h0 : _GEN_849;
  assign _GEN_851 = 10'h353 == index ? 32'h0 : _GEN_850;
  assign _GEN_852 = 10'h354 == index ? 32'h0 : _GEN_851;
  assign _GEN_853 = 10'h355 == index ? 32'h0 : _GEN_852;
  assign _GEN_854 = 10'h356 == index ? 32'h0 : _GEN_853;
  assign _GEN_855 = 10'h357 == index ? 32'h0 : _GEN_854;
  assign _GEN_856 = 10'h358 == index ? 32'h0 : _GEN_855;
  assign _GEN_857 = 10'h359 == index ? 32'h0 : _GEN_856;
  assign _GEN_858 = 10'h35a == index ? 32'h0 : _GEN_857;
  assign _GEN_859 = 10'h35b == index ? 32'h0 : _GEN_858;
  assign _GEN_860 = 10'h35c == index ? 32'h0 : _GEN_859;
  assign _GEN_861 = 10'h35d == index ? 32'h0 : _GEN_860;
  assign _GEN_862 = 10'h35e == index ? 32'h0 : _GEN_861;
  assign _GEN_863 = 10'h35f == index ? 32'h0 : _GEN_862;
  assign _GEN_864 = 10'h360 == index ? 32'h0 : _GEN_863;
  assign _GEN_865 = 10'h361 == index ? 32'h0 : _GEN_864;
  assign _GEN_866 = 10'h362 == index ? 32'h0 : _GEN_865;
  assign _GEN_867 = 10'h363 == index ? 32'h0 : _GEN_866;
  assign _GEN_868 = 10'h364 == index ? 32'h0 : _GEN_867;
  assign _GEN_869 = 10'h365 == index ? 32'h0 : _GEN_868;
  assign _GEN_870 = 10'h366 == index ? 32'h0 : _GEN_869;
  assign _GEN_871 = 10'h367 == index ? 32'h0 : _GEN_870;
  assign _GEN_872 = 10'h368 == index ? 32'h0 : _GEN_871;
  assign _GEN_873 = 10'h369 == index ? 32'h0 : _GEN_872;
  assign _GEN_874 = 10'h36a == index ? 32'h0 : _GEN_873;
  assign _GEN_875 = 10'h36b == index ? 32'h0 : _GEN_874;
  assign _GEN_876 = 10'h36c == index ? 32'h0 : _GEN_875;
  assign _GEN_877 = 10'h36d == index ? 32'h0 : _GEN_876;
  assign _GEN_878 = 10'h36e == index ? 32'h0 : _GEN_877;
  assign _GEN_879 = 10'h36f == index ? 32'h0 : _GEN_878;
  assign _GEN_880 = 10'h370 == index ? 32'h0 : _GEN_879;
  assign _GEN_881 = 10'h371 == index ? 32'h0 : _GEN_880;
  assign _GEN_882 = 10'h372 == index ? 32'h0 : _GEN_881;
  assign _GEN_883 = 10'h373 == index ? 32'h0 : _GEN_882;
  assign _GEN_884 = 10'h374 == index ? 32'h0 : _GEN_883;
  assign _GEN_885 = 10'h375 == index ? 32'h0 : _GEN_884;
  assign _GEN_886 = 10'h376 == index ? 32'h0 : _GEN_885;
  assign _GEN_887 = 10'h377 == index ? 32'h0 : _GEN_886;
  assign _GEN_888 = 10'h378 == index ? 32'h0 : _GEN_887;
  assign _GEN_889 = 10'h379 == index ? 32'h0 : _GEN_888;
  assign _GEN_890 = 10'h37a == index ? 32'h0 : _GEN_889;
  assign _GEN_891 = 10'h37b == index ? 32'h0 : _GEN_890;
  assign _GEN_892 = 10'h37c == index ? 32'h0 : _GEN_891;
  assign _GEN_893 = 10'h37d == index ? 32'h0 : _GEN_892;
  assign _GEN_894 = 10'h37e == index ? 32'h0 : _GEN_893;
  assign _GEN_895 = 10'h37f == index ? 32'h0 : _GEN_894;
  assign _GEN_896 = 10'h380 == index ? 32'h0 : _GEN_895;
  assign _GEN_897 = 10'h381 == index ? 32'h0 : _GEN_896;
  assign _GEN_898 = 10'h382 == index ? 32'h0 : _GEN_897;
  assign _GEN_899 = 10'h383 == index ? 32'h0 : _GEN_898;
  assign _GEN_900 = 10'h384 == index ? 32'h0 : _GEN_899;
  assign _GEN_901 = 10'h385 == index ? 32'h0 : _GEN_900;
  assign _GEN_902 = 10'h386 == index ? 32'h0 : _GEN_901;
  assign _GEN_903 = 10'h387 == index ? 32'h0 : _GEN_902;
  assign _GEN_904 = 10'h388 == index ? 32'h0 : _GEN_903;
  assign _GEN_905 = 10'h389 == index ? 32'h0 : _GEN_904;
  assign _GEN_906 = 10'h38a == index ? 32'h0 : _GEN_905;
  assign _GEN_907 = 10'h38b == index ? 32'h0 : _GEN_906;
  assign _GEN_908 = 10'h38c == index ? 32'h0 : _GEN_907;
  assign _GEN_909 = 10'h38d == index ? 32'h0 : _GEN_908;
  assign _GEN_910 = 10'h38e == index ? 32'h0 : _GEN_909;
  assign _GEN_911 = 10'h38f == index ? 32'h0 : _GEN_910;
  assign _GEN_912 = 10'h390 == index ? 32'h0 : _GEN_911;
  assign _GEN_913 = 10'h391 == index ? 32'h0 : _GEN_912;
  assign _GEN_914 = 10'h392 == index ? 32'h0 : _GEN_913;
  assign _GEN_915 = 10'h393 == index ? 32'h0 : _GEN_914;
  assign _GEN_916 = 10'h394 == index ? 32'h0 : _GEN_915;
  assign _GEN_917 = 10'h395 == index ? 32'h0 : _GEN_916;
  assign _GEN_918 = 10'h396 == index ? 32'h0 : _GEN_917;
  assign _GEN_919 = 10'h397 == index ? 32'h0 : _GEN_918;
  assign _GEN_920 = 10'h398 == index ? 32'h0 : _GEN_919;
  assign _GEN_921 = 10'h399 == index ? 32'h0 : _GEN_920;
  assign _GEN_922 = 10'h39a == index ? 32'h0 : _GEN_921;
  assign _GEN_923 = 10'h39b == index ? 32'h0 : _GEN_922;
  assign _GEN_924 = 10'h39c == index ? 32'h0 : _GEN_923;
  assign _GEN_925 = 10'h39d == index ? 32'h0 : _GEN_924;
  assign _GEN_926 = 10'h39e == index ? 32'h0 : _GEN_925;
  assign _GEN_927 = 10'h39f == index ? 32'h0 : _GEN_926;
  assign _GEN_928 = 10'h3a0 == index ? 32'h0 : _GEN_927;
  assign _GEN_929 = 10'h3a1 == index ? 32'h0 : _GEN_928;
  assign _GEN_930 = 10'h3a2 == index ? 32'h0 : _GEN_929;
  assign _GEN_931 = 10'h3a3 == index ? 32'h0 : _GEN_930;
  assign _GEN_932 = 10'h3a4 == index ? 32'h0 : _GEN_931;
  assign _GEN_933 = 10'h3a5 == index ? 32'h0 : _GEN_932;
  assign _GEN_934 = 10'h3a6 == index ? 32'h0 : _GEN_933;
  assign _GEN_935 = 10'h3a7 == index ? 32'h0 : _GEN_934;
  assign _GEN_936 = 10'h3a8 == index ? 32'h0 : _GEN_935;
  assign _GEN_937 = 10'h3a9 == index ? 32'h0 : _GEN_936;
  assign _GEN_938 = 10'h3aa == index ? 32'h0 : _GEN_937;
  assign _GEN_939 = 10'h3ab == index ? 32'h0 : _GEN_938;
  assign _GEN_940 = 10'h3ac == index ? 32'h0 : _GEN_939;
  assign _GEN_941 = 10'h3ad == index ? 32'h0 : _GEN_940;
  assign _GEN_942 = 10'h3ae == index ? 32'h0 : _GEN_941;
  assign _GEN_943 = 10'h3af == index ? 32'h0 : _GEN_942;
  assign _GEN_944 = 10'h3b0 == index ? 32'h0 : _GEN_943;
  assign _GEN_945 = 10'h3b1 == index ? 32'h0 : _GEN_944;
  assign _GEN_946 = 10'h3b2 == index ? 32'h0 : _GEN_945;
  assign _GEN_947 = 10'h3b3 == index ? 32'h0 : _GEN_946;
  assign _GEN_948 = 10'h3b4 == index ? 32'h0 : _GEN_947;
  assign _GEN_949 = 10'h3b5 == index ? 32'h0 : _GEN_948;
  assign _GEN_950 = 10'h3b6 == index ? 32'h0 : _GEN_949;
  assign _GEN_951 = 10'h3b7 == index ? 32'h0 : _GEN_950;
  assign _GEN_952 = 10'h3b8 == index ? 32'h0 : _GEN_951;
  assign _GEN_953 = 10'h3b9 == index ? 32'h0 : _GEN_952;
  assign _GEN_954 = 10'h3ba == index ? 32'h0 : _GEN_953;
  assign _GEN_955 = 10'h3bb == index ? 32'h0 : _GEN_954;
  assign _GEN_956 = 10'h3bc == index ? 32'h0 : _GEN_955;
  assign _GEN_957 = 10'h3bd == index ? 32'h0 : _GEN_956;
  assign _GEN_958 = 10'h3be == index ? 32'h0 : _GEN_957;
  assign _GEN_959 = 10'h3bf == index ? 32'h0 : _GEN_958;
  assign _GEN_960 = 10'h3c0 == index ? 32'h0 : _GEN_959;
  assign _GEN_961 = 10'h3c1 == index ? 32'h0 : _GEN_960;
  assign _GEN_962 = 10'h3c2 == index ? 32'h0 : _GEN_961;
  assign _GEN_963 = 10'h3c3 == index ? 32'h0 : _GEN_962;
  assign _GEN_964 = 10'h3c4 == index ? 32'h0 : _GEN_963;
  assign _GEN_965 = 10'h3c5 == index ? 32'h0 : _GEN_964;
  assign _GEN_966 = 10'h3c6 == index ? 32'h0 : _GEN_965;
  assign _GEN_967 = 10'h3c7 == index ? 32'h0 : _GEN_966;
  assign _GEN_968 = 10'h3c8 == index ? 32'h0 : _GEN_967;
  assign _GEN_969 = 10'h3c9 == index ? 32'h0 : _GEN_968;
  assign _GEN_970 = 10'h3ca == index ? 32'h0 : _GEN_969;
  assign _GEN_971 = 10'h3cb == index ? 32'h0 : _GEN_970;
  assign _GEN_972 = 10'h3cc == index ? 32'h0 : _GEN_971;
  assign _GEN_973 = 10'h3cd == index ? 32'h0 : _GEN_972;
  assign _GEN_974 = 10'h3ce == index ? 32'h0 : _GEN_973;
  assign _GEN_975 = 10'h3cf == index ? 32'h0 : _GEN_974;
  assign _GEN_976 = 10'h3d0 == index ? 32'h0 : _GEN_975;
  assign _GEN_977 = 10'h3d1 == index ? 32'h0 : _GEN_976;
  assign _GEN_978 = 10'h3d2 == index ? 32'h0 : _GEN_977;
  assign _GEN_979 = 10'h3d3 == index ? 32'h0 : _GEN_978;
  assign _GEN_980 = 10'h3d4 == index ? 32'h0 : _GEN_979;
  assign _GEN_981 = 10'h3d5 == index ? 32'h0 : _GEN_980;
  assign _GEN_982 = 10'h3d6 == index ? 32'h0 : _GEN_981;
  assign _GEN_983 = 10'h3d7 == index ? 32'h0 : _GEN_982;
  assign _GEN_984 = 10'h3d8 == index ? 32'h0 : _GEN_983;
  assign _GEN_985 = 10'h3d9 == index ? 32'h0 : _GEN_984;
  assign _GEN_986 = 10'h3da == index ? 32'h0 : _GEN_985;
  assign _GEN_987 = 10'h3db == index ? 32'h0 : _GEN_986;
  assign _GEN_988 = 10'h3dc == index ? 32'h0 : _GEN_987;
  assign _GEN_989 = 10'h3dd == index ? 32'h0 : _GEN_988;
  assign _GEN_990 = 10'h3de == index ? 32'h0 : _GEN_989;
  assign _GEN_991 = 10'h3df == index ? 32'h0 : _GEN_990;
  assign _GEN_992 = 10'h3e0 == index ? 32'h0 : _GEN_991;
  assign _GEN_993 = 10'h3e1 == index ? 32'h0 : _GEN_992;
  assign _GEN_994 = 10'h3e2 == index ? 32'h0 : _GEN_993;
  assign _GEN_995 = 10'h3e3 == index ? 32'h0 : _GEN_994;
  assign _GEN_996 = 10'h3e4 == index ? 32'h0 : _GEN_995;
  assign _GEN_997 = 10'h3e5 == index ? 32'h0 : _GEN_996;
  assign _GEN_998 = 10'h3e6 == index ? 32'h0 : _GEN_997;
  assign _GEN_999 = 10'h3e7 == index ? 32'h0 : _GEN_998;
  assign _GEN_1000 = 10'h3e8 == index ? 32'h0 : _GEN_999;
  assign _GEN_1001 = 10'h3e9 == index ? 32'h0 : _GEN_1000;
  assign _GEN_1002 = 10'h3ea == index ? 32'h0 : _GEN_1001;
  assign _GEN_1003 = 10'h3eb == index ? 32'h0 : _GEN_1002;
  assign _GEN_1004 = 10'h3ec == index ? 32'h0 : _GEN_1003;
  assign _GEN_1005 = 10'h3ed == index ? 32'h0 : _GEN_1004;
  assign _GEN_1006 = 10'h3ee == index ? 32'h0 : _GEN_1005;
  assign _GEN_1007 = 10'h3ef == index ? 32'h0 : _GEN_1006;
  assign _GEN_1008 = 10'h3f0 == index ? 32'h0 : _GEN_1007;
  assign _GEN_1009 = 10'h3f1 == index ? 32'h0 : _GEN_1008;
  assign _GEN_1010 = 10'h3f2 == index ? 32'h0 : _GEN_1009;
  assign _GEN_1011 = 10'h3f3 == index ? 32'h0 : _GEN_1010;
  assign _GEN_1012 = 10'h3f4 == index ? 32'h0 : _GEN_1011;
  assign _GEN_1013 = 10'h3f5 == index ? 32'h0 : _GEN_1012;
  assign _GEN_1014 = 10'h3f6 == index ? 32'h0 : _GEN_1013;
  assign _GEN_1015 = 10'h3f7 == index ? 32'h0 : _GEN_1014;
  assign _GEN_1016 = 10'h3f8 == index ? 32'h0 : _GEN_1015;
  assign _GEN_1017 = 10'h3f9 == index ? 32'h0 : _GEN_1016;
  assign _GEN_1018 = 10'h3fa == index ? 32'h0 : _GEN_1017;
  assign _GEN_1019 = 10'h3fb == index ? 32'h0 : _GEN_1018;
  assign _GEN_1020 = 10'h3fc == index ? 32'h0 : _GEN_1019;
  assign _GEN_1021 = 10'h3fd == index ? 32'h0 : _GEN_1020;
  assign _GEN_1022 = 10'h3fe == index ? 32'h0 : _GEN_1021;
  assign _GEN_1023 = 10'h3ff == index ? 32'h0 : _GEN_1022;
  assign _T_2116 = _T_2113 ? 32'h0 : _GEN_1023;
endmodule
module Queue_41(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [3:0] io_enq_bits_size,
  input  [4:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_2;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _T_31;
  assign io_deq_bits_opcode = ram_opcode__T_35_data;
  assign io_deq_bits_size = ram_size__T_35_data;
  assign io_deq_bits_source = ram_source__T_35_data;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _T_21;
  assign ram_opcode__T_26_en = _T_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _T_21;
  assign ram_size__T_26_en = _T_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _T_21;
  assign ram_source__T_26_en = _T_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _T_21 != _T_23;
  assign _GEN_10 = _T_29 ? _T_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        maybe_full <= _T_21;
      end
    end
  end
endmodule
module Queue_42(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_param,
  input  [3:0] io_enq_bits_size,
  input  [4:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_param,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source
);
  reg [2:0] ram_param [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_param__T_35_data;
  wire  ram_param__T_35_addr;
  wire [2:0] ram_param__T_26_data;
  wire  ram_param__T_26_addr;
  wire  ram_param__T_26_mask;
  wire  ram_param__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_2;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _T_31;
  assign io_deq_bits_param = ram_param__T_35_data;
  assign io_deq_bits_size = ram_size__T_35_data;
  assign io_deq_bits_source = ram_source__T_35_data;
  assign ram_param__T_35_addr = 1'h0;
  assign ram_param__T_35_data = ram_param[ram_param__T_35_addr];
  assign ram_param__T_26_data = io_enq_bits_param;
  assign ram_param__T_26_addr = 1'h0;
  assign ram_param__T_26_mask = _T_21;
  assign ram_param__T_26_en = _T_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _T_21;
  assign ram_size__T_26_en = _T_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _T_21;
  assign ram_source__T_26_en = _T_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _T_21 != _T_23;
  assign _GEN_10 = _T_29 ? _T_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_param__T_26_en & ram_param__T_26_mask) begin
      ram_param[ram_param__T_26_addr] <= ram_param__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        maybe_full <= _T_21;
      end
    end
  end
endmodule
module TLError_error(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [3:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input         io_in_0_c_valid,
  input  [2:0]  io_in_0_c_bits_param,
  input  [3:0]  io_in_0_c_bits_size,
  input  [4:0]  io_in_0_c_bits_source,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [3:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error
);
  wire  a_clock;
  wire  a_reset;
  wire  a_io_enq_ready;
  wire  a_io_enq_valid;
  wire [2:0] a_io_enq_bits_opcode;
  wire [3:0] a_io_enq_bits_size;
  wire [4:0] a_io_enq_bits_source;
  wire  a_io_deq_ready;
  wire  a_io_deq_valid;
  wire [2:0] a_io_deq_bits_opcode;
  wire [3:0] a_io_deq_bits_size;
  wire [4:0] a_io_deq_bits_source;
  wire  c_clock;
  wire  c_reset;
  wire  c_io_enq_ready;
  wire  c_io_enq_valid;
  wire [2:0] c_io_enq_bits_param;
  wire [3:0] c_io_enq_bits_size;
  wire [4:0] c_io_enq_bits_source;
  wire  c_io_deq_ready;
  wire  c_io_deq_valid;
  wire [2:0] c_io_deq_bits_param;
  wire [3:0] c_io_deq_bits_size;
  wire [4:0] c_io_deq_bits_source;
  wire [3:0] da_bits_size;
  wire [4:0] da_bits_source;
  wire [3:0] dc_bits_size;
  wire [4:0] dc_bits_source;
  wire  _T_68;
  wire [26:0] _T_71;
  wire [11:0] _T_72;
  wire [11:0] _T_73;
  wire [9:0] _T_74;
  wire  _T_75;
  wire  _T_77;
  wire [9:0] _T_79;
  reg [9:0] _T_82;
  reg [31:0] _RAND_0;
  wire [10:0] _T_84;
  wire [10:0] _T_85;
  wire [9:0] _T_86;
  wire  _T_88;
  wire  _T_90;
  wire  _T_92;
  wire  a_last;
  wire [9:0] _T_96;
  wire [9:0] _GEN_2;
  wire  _T_125;
  wire [26:0] _T_128;
  wire [11:0] _T_129;
  wire [11:0] _T_130;
  wire [9:0] _T_131;
  wire  _T_132;
  wire [9:0] _T_134;
  reg [9:0] _T_137;
  reg [31:0] _RAND_1;
  wire [10:0] _T_139;
  wire [10:0] _T_140;
  wire [9:0] _T_141;
  wire  _T_143;
  wire  _T_145;
  wire  _T_147;
  wire  da_last;
  wire [9:0] _T_151;
  wire [9:0] _GEN_4;
  wire  _T_179;
  wire  _T_181;
  wire  _T_182;
  wire  _T_183;
  wire [2:0] _GEN_7;
  wire [2:0] _GEN_8;
  wire [2:0] _GEN_9;
  wire [2:0] _GEN_10;
  wire [2:0] _GEN_11;
  wire  _T_211;
  wire [1:0] _T_225;
  wire [1:0] _GEN_13;
  reg [9:0] _T_249;
  reg [31:0] _RAND_2;
  wire  _T_251;
  wire  _T_252;
  wire [1:0] _T_253;
  wire [2:0] _GEN_14;
  wire [2:0] _T_254;
  wire [1:0] _T_255;
  wire [1:0] _T_256;
  wire [2:0] _GEN_15;
  wire [2:0] _T_258;
  wire [1:0] _T_259;
  wire [1:0] _T_260;
  wire  _T_261;
  wire  _T_262;
  wire  _T_270;
  wire  _T_271;
  wire  _T_281;
  wire  _T_285;
  wire  _T_290;
  wire  _T_291;
  wire  _T_293;
  wire  _T_295;
  wire  _T_296;
  wire  _T_298;
  wire  _T_300;
  wire  _T_301;
  wire  _T_303;
  wire [9:0] _T_307;
  wire  _T_309;
  wire [9:0] _GEN_16;
  wire [10:0] _T_310;
  wire [10:0] _T_311;
  wire [9:0] _T_312;
  wire [9:0] _T_313;
  reg  _T_331_0;
  reg [31:0] _RAND_3;
  reg  _T_331_1;
  reg [31:0] _RAND_4;
  wire  _T_342_0;
  wire  _T_342_1;
  wire  _T_350_0;
  wire  _T_350_1;
  wire  _T_358;
  wire  _T_359;
  wire  _T_363;
  wire  _T_365;
  wire  _T_366;
  wire  _T_369;
  wire [8:0] _T_373;
  wire [4:0] _T_374;
  wire [13:0] _T_375;
  wire [47:0] _T_376;
  wire [47:0] _T_378;
  wire [8:0] _T_381;
  wire [4:0] _T_382;
  wire [13:0] _T_383;
  wire [47:0] _T_384;
  wire [47:0] _T_386;
  wire [47:0] _T_387;
  wire  _T_392;
  wire [31:0] _T_393;
  wire  _T_394;
  wire [4:0] _T_395;
  wire [3:0] _T_396;
  wire [1:0] _T_397;
  wire [2:0] _T_398;
  Queue_41 a (
    .clock(a_clock),
    .reset(a_reset),
    .io_enq_ready(a_io_enq_ready),
    .io_enq_valid(a_io_enq_valid),
    .io_enq_bits_opcode(a_io_enq_bits_opcode),
    .io_enq_bits_size(a_io_enq_bits_size),
    .io_enq_bits_source(a_io_enq_bits_source),
    .io_deq_ready(a_io_deq_ready),
    .io_deq_valid(a_io_deq_valid),
    .io_deq_bits_opcode(a_io_deq_bits_opcode),
    .io_deq_bits_size(a_io_deq_bits_size),
    .io_deq_bits_source(a_io_deq_bits_source)
  );
  Queue_42 c (
    .clock(c_clock),
    .reset(c_reset),
    .io_enq_ready(c_io_enq_ready),
    .io_enq_valid(c_io_enq_valid),
    .io_enq_bits_param(c_io_enq_bits_param),
    .io_enq_bits_size(c_io_enq_bits_size),
    .io_enq_bits_source(c_io_enq_bits_source),
    .io_deq_ready(c_io_deq_ready),
    .io_deq_valid(c_io_deq_valid),
    .io_deq_bits_param(c_io_deq_bits_param),
    .io_deq_bits_size(c_io_deq_bits_size),
    .io_deq_bits_source(c_io_deq_bits_source)
  );
  assign io_in_0_a_ready = a_io_enq_ready;
  assign io_in_0_d_valid = _T_369;
  assign io_in_0_d_bits_opcode = _T_398;
  assign io_in_0_d_bits_param = _T_397;
  assign io_in_0_d_bits_size = _T_396;
  assign io_in_0_d_bits_source = _T_395;
  assign io_in_0_d_bits_sink = _T_394;
  assign io_in_0_d_bits_data = _T_393;
  assign io_in_0_d_bits_error = _T_392;
  assign a_clock = clock;
  assign a_reset = reset;
  assign a_io_enq_valid = io_in_0_a_valid;
  assign a_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign a_io_enq_bits_size = io_in_0_a_bits_size;
  assign a_io_enq_bits_source = io_in_0_a_bits_source;
  assign a_io_deq_ready = _T_182;
  assign c_clock = clock;
  assign c_reset = reset;
  assign c_io_enq_valid = io_in_0_c_valid;
  assign c_io_enq_bits_param = io_in_0_c_bits_param;
  assign c_io_enq_bits_size = io_in_0_c_bits_size;
  assign c_io_enq_bits_source = io_in_0_c_bits_source;
  assign c_io_deq_ready = _T_358;
  assign da_bits_size = a_io_deq_bits_size;
  assign da_bits_source = a_io_deq_bits_source;
  assign dc_bits_size = c_io_deq_bits_size;
  assign dc_bits_source = c_io_deq_bits_source;
  assign _T_68 = a_io_deq_ready & a_io_deq_valid;
  assign _T_71 = 27'hfff << a_io_deq_bits_size;
  assign _T_72 = _T_71[11:0];
  assign _T_73 = ~ _T_72;
  assign _T_74 = _T_73[11:2];
  assign _T_75 = a_io_deq_bits_opcode[2];
  assign _T_77 = _T_75 == 1'h0;
  assign _T_79 = _T_77 ? _T_74 : 10'h0;
  assign _T_84 = _T_82 - 10'h1;
  assign _T_85 = $unsigned(_T_84);
  assign _T_86 = _T_85[9:0];
  assign _T_88 = _T_82 == 10'h0;
  assign _T_90 = _T_82 == 10'h1;
  assign _T_92 = _T_79 == 10'h0;
  assign a_last = _T_90 | _T_92;
  assign _T_96 = _T_88 ? _T_79 : _T_86;
  assign _GEN_2 = _T_68 ? _T_96 : _T_82;
  assign _T_125 = _T_359 & _T_183;
  assign _T_128 = 27'hfff << da_bits_size;
  assign _T_129 = _T_128[11:0];
  assign _T_130 = ~ _T_129;
  assign _T_131 = _T_130[11:2];
  assign _T_132 = _GEN_11[0];
  assign _T_134 = _T_132 ? _T_131 : 10'h0;
  assign _T_139 = _T_137 - 10'h1;
  assign _T_140 = $unsigned(_T_139);
  assign _T_141 = _T_140[9:0];
  assign _T_143 = _T_137 == 10'h0;
  assign _T_145 = _T_137 == 10'h1;
  assign _T_147 = _T_134 == 10'h0;
  assign da_last = _T_145 | _T_147;
  assign _T_151 = _T_143 ? _T_134 : _T_141;
  assign _GEN_4 = _T_125 ? _T_151 : _T_137;
  assign _T_179 = _T_359 & da_last;
  assign _T_181 = a_last == 1'h0;
  assign _T_182 = _T_179 | _T_181;
  assign _T_183 = a_io_deq_valid & a_last;
  assign _GEN_7 = 3'h2 == a_io_deq_bits_opcode ? 3'h1 : 3'h0;
  assign _GEN_8 = 3'h3 == a_io_deq_bits_opcode ? 3'h1 : _GEN_7;
  assign _GEN_9 = 3'h4 == a_io_deq_bits_opcode ? 3'h1 : _GEN_8;
  assign _GEN_10 = 3'h5 == a_io_deq_bits_opcode ? 3'h2 : _GEN_9;
  assign _GEN_11 = 3'h6 == a_io_deq_bits_opcode ? 3'h4 : _GEN_10;
  assign _T_211 = c_io_deq_valid;
  assign _T_225 = c_io_deq_bits_param[1:0];
  assign _GEN_13 = 2'h2 == _T_225 ? 2'h1 : 2'h2;
  assign _T_251 = _T_249 == 10'h0;
  assign _T_252 = _T_251 & io_in_0_d_ready;
  assign _T_253 = {_T_183,_T_211};
  assign _GEN_14 = {{1'd0}, _T_253};
  assign _T_254 = _GEN_14 << 1;
  assign _T_255 = _T_254[1:0];
  assign _T_256 = _T_253 | _T_255;
  assign _GEN_15 = {{1'd0}, _T_256};
  assign _T_258 = _GEN_15 << 1;
  assign _T_259 = _T_258[1:0];
  assign _T_260 = ~ _T_259;
  assign _T_261 = _T_260[0];
  assign _T_262 = _T_260[1];
  assign _T_270 = _T_261 & _T_211;
  assign _T_271 = _T_262 & _T_183;
  assign _T_281 = _T_270 | _T_271;
  assign _T_285 = _T_270 == 1'h0;
  assign _T_290 = _T_271 == 1'h0;
  assign _T_291 = _T_285 | _T_290;
  assign _T_293 = _T_291 | reset;
  assign _T_295 = _T_293 == 1'h0;
  assign _T_296 = _T_211 | _T_183;
  assign _T_298 = _T_296 == 1'h0;
  assign _T_300 = _T_298 | _T_281;
  assign _T_301 = _T_300 | reset;
  assign _T_303 = _T_301 == 1'h0;
  assign _T_307 = _T_271 ? _T_134 : 10'h0;
  assign _T_309 = io_in_0_d_ready & io_in_0_d_valid;
  assign _GEN_16 = {{9'd0}, _T_309};
  assign _T_310 = _T_249 - _GEN_16;
  assign _T_311 = $unsigned(_T_310);
  assign _T_312 = _T_311[9:0];
  assign _T_313 = _T_252 ? _T_307 : _T_312;
  assign _T_342_0 = _T_251 ? _T_270 : _T_331_0;
  assign _T_342_1 = _T_251 ? _T_271 : _T_331_1;
  assign _T_350_0 = _T_251 ? _T_261 : _T_331_0;
  assign _T_350_1 = _T_251 ? _T_262 : _T_331_1;
  assign _T_358 = io_in_0_d_ready & _T_350_0;
  assign _T_359 = io_in_0_d_ready & _T_350_1;
  assign _T_363 = _T_331_0 ? _T_211 : 1'h0;
  assign _T_365 = _T_331_1 ? _T_183 : 1'h0;
  assign _T_366 = _T_363 | _T_365;
  assign _T_369 = _T_251 ? _T_296 : _T_366;
  assign _T_373 = {dc_bits_size,dc_bits_source};
  assign _T_374 = {3'h6,_GEN_13};
  assign _T_375 = {_T_374,_T_373};
  assign _T_376 = {_T_375,34'h1};
  assign _T_378 = _T_342_0 ? _T_376 : 48'h0;
  assign _T_381 = {da_bits_size,da_bits_source};
  assign _T_382 = {_GEN_11,2'h0};
  assign _T_383 = {_T_382,_T_381};
  assign _T_384 = {_T_383,34'h1};
  assign _T_386 = _T_342_1 ? _T_384 : 48'h0;
  assign _T_387 = _T_378 | _T_386;
  assign _T_392 = _T_387[0];
  assign _T_393 = _T_387[32:1];
  assign _T_394 = _T_387[33];
  assign _T_395 = _T_387[38:34];
  assign _T_396 = _T_387[42:39];
  assign _T_397 = _T_387[44:43];
  assign _T_398 = _T_387[47:45];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_82 = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_137 = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_249 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_331_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_331_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_82 <= 10'h0;
    end else begin
      if (_T_68) begin
        if (_T_88) begin
          if (_T_77) begin
            _T_82 <= _T_74;
          end else begin
            _T_82 <= 10'h0;
          end
        end else begin
          _T_82 <= _T_86;
        end
      end
    end
    if (reset) begin
      _T_137 <= 10'h0;
    end else begin
      if (_T_125) begin
        if (_T_143) begin
          if (_T_132) begin
            _T_137 <= _T_131;
          end else begin
            _T_137 <= 10'h0;
          end
        end else begin
          _T_137 <= _T_141;
        end
      end
    end
    if (reset) begin
      _T_249 <= 10'h0;
    end else begin
      if (_T_252) begin
        if (_T_271) begin
          if (_T_132) begin
            _T_249 <= _T_131;
          end else begin
            _T_249 <= 10'h0;
          end
        end else begin
          _T_249 <= 10'h0;
        end
      end else begin
        _T_249 <= _T_312;
      end
    end
    if (reset) begin
      _T_331_0 <= 1'h0;
    end else begin
      if (_T_251) begin
        _T_331_0 <= _T_270;
      end
    end
    if (reset) begin
      _T_331_1 <= 1'h0;
    end else begin
      if (_T_251) begin
        _T_331_1 <= _T_271;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_295) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:66 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_295) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_303) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Arbiter.scala:68 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_303) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_43(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [2:0] io_enq_bits_opcode,
  input  [3:0] io_enq_bits_size,
  input  [4:0] io_enq_bits_source,
  input        io_deq_ready,
  output       io_deq_valid,
  output [2:0] io_deq_bits_opcode,
  output [3:0] io_deq_bits_size,
  output [4:0] io_deq_bits_source
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_1;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_2;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_3;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  assign io_enq_ready = _GEN_11;
  assign io_deq_valid = _T_31;
  assign io_deq_bits_opcode = ram_opcode__T_35_data;
  assign io_deq_bits_size = ram_size__T_35_data;
  assign io_deq_bits_source = ram_source__T_35_data;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _T_21;
  assign ram_opcode__T_26_en = _T_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _T_21;
  assign ram_size__T_26_en = _T_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _T_21;
  assign ram_source__T_26_en = _T_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _T_21 != _T_23;
  assign _GEN_10 = _T_29 ? _T_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_deq_ready ? 1'h1 : _T_18;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_1[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  maybe_full = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        maybe_full <= _T_21;
      end
    end
  end
endmodule
module Queue_44(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [2:0]  io_enq_bits_opcode,
  input  [1:0]  io_enq_bits_param,
  input  [3:0]  io_enq_bits_size,
  input  [4:0]  io_enq_bits_source,
  input         io_enq_bits_sink,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_error,
  input         io_deq_ready,
  output        io_deq_valid,
  output [2:0]  io_deq_bits_opcode,
  output [1:0]  io_deq_bits_param,
  output [3:0]  io_deq_bits_size,
  output [4:0]  io_deq_bits_source,
  output        io_deq_bits_sink,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_error
);
  reg [2:0] ram_opcode [0:0];
  reg [31:0] _RAND_0;
  wire [2:0] ram_opcode__T_35_data;
  wire  ram_opcode__T_35_addr;
  wire [2:0] ram_opcode__T_26_data;
  wire  ram_opcode__T_26_addr;
  wire  ram_opcode__T_26_mask;
  wire  ram_opcode__T_26_en;
  reg [1:0] ram_param [0:0];
  reg [31:0] _RAND_1;
  wire [1:0] ram_param__T_35_data;
  wire  ram_param__T_35_addr;
  wire [1:0] ram_param__T_26_data;
  wire  ram_param__T_26_addr;
  wire  ram_param__T_26_mask;
  wire  ram_param__T_26_en;
  reg [3:0] ram_size [0:0];
  reg [31:0] _RAND_2;
  wire [3:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [3:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [4:0] ram_source [0:0];
  reg [31:0] _RAND_3;
  wire [4:0] ram_source__T_35_data;
  wire  ram_source__T_35_addr;
  wire [4:0] ram_source__T_26_data;
  wire  ram_source__T_26_addr;
  wire  ram_source__T_26_mask;
  wire  ram_source__T_26_en;
  reg  ram_sink [0:0];
  reg [31:0] _RAND_4;
  wire  ram_sink__T_35_data;
  wire  ram_sink__T_35_addr;
  wire  ram_sink__T_26_data;
  wire  ram_sink__T_26_addr;
  wire  ram_sink__T_26_mask;
  wire  ram_sink__T_26_en;
  reg [31:0] ram_data [0:0];
  reg [31:0] _RAND_5;
  wire [31:0] ram_data__T_35_data;
  wire  ram_data__T_35_addr;
  wire [31:0] ram_data__T_26_data;
  wire  ram_data__T_26_addr;
  wire  ram_data__T_26_mask;
  wire  ram_data__T_26_en;
  reg  ram_error [0:0];
  reg [31:0] _RAND_6;
  wire  ram_error__T_35_data;
  wire  ram_error__T_35_addr;
  wire  ram_error__T_26_data;
  wire  ram_error__T_26_addr;
  wire  ram_error__T_26_mask;
  wire  ram_error__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_10;
  wire  _T_31;
  wire  _GEN_11;
  assign io_enq_ready = _GEN_11;
  assign io_deq_valid = _T_31;
  assign io_deq_bits_opcode = ram_opcode__T_35_data;
  assign io_deq_bits_param = ram_param__T_35_data;
  assign io_deq_bits_size = ram_size__T_35_data;
  assign io_deq_bits_source = ram_source__T_35_data;
  assign io_deq_bits_sink = ram_sink__T_35_data;
  assign io_deq_bits_data = ram_data__T_35_data;
  assign io_deq_bits_error = ram_error__T_35_data;
  assign ram_opcode__T_35_addr = 1'h0;
  assign ram_opcode__T_35_data = ram_opcode[ram_opcode__T_35_addr];
  assign ram_opcode__T_26_data = io_enq_bits_opcode;
  assign ram_opcode__T_26_addr = 1'h0;
  assign ram_opcode__T_26_mask = _T_21;
  assign ram_opcode__T_26_en = _T_21;
  assign ram_param__T_35_addr = 1'h0;
  assign ram_param__T_35_data = ram_param[ram_param__T_35_addr];
  assign ram_param__T_26_data = io_enq_bits_param;
  assign ram_param__T_26_addr = 1'h0;
  assign ram_param__T_26_mask = _T_21;
  assign ram_param__T_26_en = _T_21;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _T_21;
  assign ram_size__T_26_en = _T_21;
  assign ram_source__T_35_addr = 1'h0;
  assign ram_source__T_35_data = ram_source[ram_source__T_35_addr];
  assign ram_source__T_26_data = io_enq_bits_source;
  assign ram_source__T_26_addr = 1'h0;
  assign ram_source__T_26_mask = _T_21;
  assign ram_source__T_26_en = _T_21;
  assign ram_sink__T_35_addr = 1'h0;
  assign ram_sink__T_35_data = ram_sink[ram_sink__T_35_addr];
  assign ram_sink__T_26_data = io_enq_bits_sink;
  assign ram_sink__T_26_addr = 1'h0;
  assign ram_sink__T_26_mask = _T_21;
  assign ram_sink__T_26_en = _T_21;
  assign ram_data__T_35_addr = 1'h0;
  assign ram_data__T_35_data = ram_data[ram_data__T_35_addr];
  assign ram_data__T_26_data = io_enq_bits_data;
  assign ram_data__T_26_addr = 1'h0;
  assign ram_data__T_26_mask = _T_21;
  assign ram_data__T_26_en = _T_21;
  assign ram_error__T_35_addr = 1'h0;
  assign ram_error__T_35_data = ram_error[ram_error__T_35_addr];
  assign ram_error__T_26_data = io_enq_bits_error;
  assign ram_error__T_26_addr = 1'h0;
  assign ram_error__T_26_mask = _T_21;
  assign ram_error__T_26_en = _T_21;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _T_21 != _T_23;
  assign _GEN_10 = _T_29 ? _T_21 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_11 = io_deq_ready ? 1'h1 : _T_18;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_opcode[initvar] = _RAND_0[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_param[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_2[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_source[initvar] = _RAND_3[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_sink[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_error[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_opcode__T_26_en & ram_opcode__T_26_mask) begin
      ram_opcode[ram_opcode__T_26_addr] <= ram_opcode__T_26_data;
    end
    if(ram_param__T_26_en & ram_param__T_26_mask) begin
      ram_param[ram_param__T_26_addr] <= ram_param__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_source__T_26_en & ram_source__T_26_mask) begin
      ram_source[ram_source__T_26_addr] <= ram_source__T_26_data;
    end
    if(ram_sink__T_26_en & ram_sink__T_26_mask) begin
      ram_sink[ram_sink__T_26_addr] <= ram_sink__T_26_data;
    end
    if(ram_data__T_26_en & ram_data__T_26_mask) begin
      ram_data[ram_data__T_26_addr] <= ram_data__T_26_data;
    end
    if(ram_error__T_26_en & ram_error__T_26_mask) begin
      ram_error[ram_error__T_26_addr] <= ram_error__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        maybe_full <= _T_21;
      end
    end
  end
endmodule
module TLBuffer_error(
  input         clock,
  input         reset,
  output        io_in_0_a_ready,
  input         io_in_0_a_valid,
  input  [2:0]  io_in_0_a_bits_opcode,
  input  [3:0]  io_in_0_a_bits_size,
  input  [4:0]  io_in_0_a_bits_source,
  input         io_in_0_d_ready,
  output        io_in_0_d_valid,
  output [2:0]  io_in_0_d_bits_opcode,
  output [1:0]  io_in_0_d_bits_param,
  output [3:0]  io_in_0_d_bits_size,
  output [4:0]  io_in_0_d_bits_source,
  output        io_in_0_d_bits_sink,
  output [31:0] io_in_0_d_bits_data,
  output        io_in_0_d_bits_error,
  input         io_out_0_a_ready,
  output        io_out_0_a_valid,
  output [2:0]  io_out_0_a_bits_opcode,
  output [3:0]  io_out_0_a_bits_size,
  output [4:0]  io_out_0_a_bits_source,
  output        io_out_0_c_valid,
  output [2:0]  io_out_0_c_bits_param,
  output [3:0]  io_out_0_c_bits_size,
  output [4:0]  io_out_0_c_bits_source,
  output        io_out_0_d_ready,
  input         io_out_0_d_valid,
  input  [2:0]  io_out_0_d_bits_opcode,
  input  [1:0]  io_out_0_d_bits_param,
  input  [3:0]  io_out_0_d_bits_size,
  input  [4:0]  io_out_0_d_bits_source,
  input         io_out_0_d_bits_sink,
  input  [31:0] io_out_0_d_bits_data,
  input         io_out_0_d_bits_error
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [2:0] Queue_io_enq_bits_opcode;
  wire [3:0] Queue_io_enq_bits_size;
  wire [4:0] Queue_io_enq_bits_source;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [2:0] Queue_io_deq_bits_opcode;
  wire [3:0] Queue_io_deq_bits_size;
  wire [4:0] Queue_io_deq_bits_source;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [2:0] Queue_1_io_enq_bits_opcode;
  wire [1:0] Queue_1_io_enq_bits_param;
  wire [3:0] Queue_1_io_enq_bits_size;
  wire [4:0] Queue_1_io_enq_bits_source;
  wire  Queue_1_io_enq_bits_sink;
  wire [31:0] Queue_1_io_enq_bits_data;
  wire  Queue_1_io_enq_bits_error;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [2:0] Queue_1_io_deq_bits_opcode;
  wire [1:0] Queue_1_io_deq_bits_param;
  wire [3:0] Queue_1_io_deq_bits_size;
  wire [4:0] Queue_1_io_deq_bits_source;
  wire  Queue_1_io_deq_bits_sink;
  wire [31:0] Queue_1_io_deq_bits_data;
  wire  Queue_1_io_deq_bits_error;
  Queue_43 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_opcode(Queue_io_enq_bits_opcode),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_source(Queue_io_enq_bits_source),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_opcode(Queue_io_deq_bits_opcode),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_source(Queue_io_deq_bits_source)
  );
  Queue_44 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_opcode(Queue_1_io_enq_bits_opcode),
    .io_enq_bits_param(Queue_1_io_enq_bits_param),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_source(Queue_1_io_enq_bits_source),
    .io_enq_bits_sink(Queue_1_io_enq_bits_sink),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_error(Queue_1_io_enq_bits_error),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_opcode(Queue_1_io_deq_bits_opcode),
    .io_deq_bits_param(Queue_1_io_deq_bits_param),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_source(Queue_1_io_deq_bits_source),
    .io_deq_bits_sink(Queue_1_io_deq_bits_sink),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_error(Queue_1_io_deq_bits_error)
  );
  assign io_in_0_a_ready = Queue_io_enq_ready;
  assign io_in_0_d_valid = Queue_1_io_deq_valid;
  assign io_in_0_d_bits_opcode = Queue_1_io_deq_bits_opcode;
  assign io_in_0_d_bits_param = Queue_1_io_deq_bits_param;
  assign io_in_0_d_bits_size = Queue_1_io_deq_bits_size;
  assign io_in_0_d_bits_source = Queue_1_io_deq_bits_source;
  assign io_in_0_d_bits_sink = Queue_1_io_deq_bits_sink;
  assign io_in_0_d_bits_data = Queue_1_io_deq_bits_data;
  assign io_in_0_d_bits_error = Queue_1_io_deq_bits_error;
  assign io_out_0_a_valid = Queue_io_deq_valid;
  assign io_out_0_a_bits_opcode = Queue_io_deq_bits_opcode;
  assign io_out_0_a_bits_size = Queue_io_deq_bits_size;
  assign io_out_0_a_bits_source = Queue_io_deq_bits_source;
  assign io_out_0_c_valid = 1'h0;
  assign io_out_0_c_bits_param = 3'h0;
  assign io_out_0_c_bits_size = 4'h0;
  assign io_out_0_c_bits_source = 5'h0;
  assign io_out_0_d_ready = Queue_1_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_a_valid;
  assign Queue_io_enq_bits_opcode = io_in_0_a_bits_opcode;
  assign Queue_io_enq_bits_size = io_in_0_a_bits_size;
  assign Queue_io_enq_bits_source = io_in_0_a_bits_source;
  assign Queue_io_deq_ready = io_out_0_a_ready;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_out_0_d_valid;
  assign Queue_1_io_enq_bits_opcode = io_out_0_d_bits_opcode;
  assign Queue_1_io_enq_bits_param = io_out_0_d_bits_param;
  assign Queue_1_io_enq_bits_size = io_out_0_d_bits_size;
  assign Queue_1_io_enq_bits_source = io_out_0_d_bits_source;
  assign Queue_1_io_enq_bits_sink = io_out_0_d_bits_sink;
  assign Queue_1_io_enq_bits_data = io_out_0_d_bits_data;
  assign Queue_1_io_enq_bits_error = io_out_0_d_bits_error;
  assign Queue_1_io_deq_ready = io_in_0_d_ready;
endmodule
module ExampleRocketSystem(
  input         clock,
  input         reset,
  output        debug_clockeddmi_dmi_req_ready,
  input         debug_clockeddmi_dmi_req_valid,
  input  [6:0]  debug_clockeddmi_dmi_req_bits_addr,
  input  [31:0] debug_clockeddmi_dmi_req_bits_data,
  input  [1:0]  debug_clockeddmi_dmi_req_bits_op,
  input         debug_clockeddmi_dmi_resp_ready,
  output        debug_clockeddmi_dmi_resp_valid,
  output [31:0] debug_clockeddmi_dmi_resp_bits_data,
  output [1:0]  debug_clockeddmi_dmi_resp_bits_resp,
  input         debug_clockeddmi_dmiClock,
  input         debug_clockeddmi_dmiReset,
  output        debug_ndreset,
  input  [1:0]  interrupts,
  input         mmio_axi4_0_aw_ready,
  output        mmio_axi4_0_aw_valid,
  output [3:0]  mmio_axi4_0_aw_bits_id,
  output [30:0] mmio_axi4_0_aw_bits_addr,
  output [7:0]  mmio_axi4_0_aw_bits_len,
  output [2:0]  mmio_axi4_0_aw_bits_size,
  output [1:0]  mmio_axi4_0_aw_bits_burst,
  input         mmio_axi4_0_w_ready,
  output        mmio_axi4_0_w_valid,
  output [63:0] mmio_axi4_0_w_bits_data,
  output [7:0]  mmio_axi4_0_w_bits_strb,
  output        mmio_axi4_0_w_bits_last,
  output        mmio_axi4_0_b_ready,
  input         mmio_axi4_0_b_valid,
  input  [3:0]  mmio_axi4_0_b_bits_id,
  input  [1:0]  mmio_axi4_0_b_bits_resp,
  input         mmio_axi4_0_ar_ready,
  output        mmio_axi4_0_ar_valid,
  output [3:0]  mmio_axi4_0_ar_bits_id,
  output [30:0] mmio_axi4_0_ar_bits_addr,
  output [7:0]  mmio_axi4_0_ar_bits_len,
  output [2:0]  mmio_axi4_0_ar_bits_size,
  output [1:0]  mmio_axi4_0_ar_bits_burst,
  output        mmio_axi4_0_r_ready,
  input         mmio_axi4_0_r_valid,
  input  [3:0]  mmio_axi4_0_r_bits_id,
  input  [63:0] mmio_axi4_0_r_bits_data,
  input  [1:0]  mmio_axi4_0_r_bits_resp,
  input         mmio_axi4_0_r_bits_last,
  input         l2_frontend_bus_axi4_0_aw_valid,
  input  [7:0]  l2_frontend_bus_axi4_0_aw_bits_id,
  input  [31:0] l2_frontend_bus_axi4_0_aw_bits_addr,
  input  [7:0]  l2_frontend_bus_axi4_0_aw_bits_len,
  input  [2:0]  l2_frontend_bus_axi4_0_aw_bits_size,
  input  [1:0]  l2_frontend_bus_axi4_0_aw_bits_burst,
  input         l2_frontend_bus_axi4_0_w_valid,
  input  [63:0] l2_frontend_bus_axi4_0_w_bits_data,
  input  [7:0]  l2_frontend_bus_axi4_0_w_bits_strb,
  input         l2_frontend_bus_axi4_0_w_bits_last,
  input         l2_frontend_bus_axi4_0_b_ready,
  input         l2_frontend_bus_axi4_0_ar_valid,
  input  [7:0]  l2_frontend_bus_axi4_0_ar_bits_id,
  input  [31:0] l2_frontend_bus_axi4_0_ar_bits_addr,
  input  [7:0]  l2_frontend_bus_axi4_0_ar_bits_len,
  input  [2:0]  l2_frontend_bus_axi4_0_ar_bits_size,
  input  [1:0]  l2_frontend_bus_axi4_0_ar_bits_burst,
  input         l2_frontend_bus_axi4_0_r_ready
);
  wire  IntXbar_io_in_0_0;
  wire  IntXbar_io_in_0_1;
  wire  IntXbar_io_out_0_0;
  wire  IntXbar_io_out_0_1;
  wire  TLXbar_clock;
  wire  TLXbar_reset;
  wire  TLXbar_io_in_1_a_ready;
  wire  TLXbar_io_in_1_a_valid;
  wire [2:0] TLXbar_io_in_1_a_bits_opcode;
  wire [2:0] TLXbar_io_in_1_a_bits_param;
  wire [3:0] TLXbar_io_in_1_a_bits_size;
  wire [3:0] TLXbar_io_in_1_a_bits_source;
  wire [31:0] TLXbar_io_in_1_a_bits_address;
  wire [3:0] TLXbar_io_in_1_a_bits_mask;
  wire [31:0] TLXbar_io_in_1_a_bits_data;
  wire  TLXbar_io_in_1_d_ready;
  wire  TLXbar_io_in_1_d_valid;
  wire [2:0] TLXbar_io_in_1_d_bits_opcode;
  wire [3:0] TLXbar_io_in_1_d_bits_size;
  wire [3:0] TLXbar_io_in_1_d_bits_source;
  wire  TLXbar_io_in_0_a_ready;
  wire  TLXbar_io_in_0_a_valid;
  wire [2:0] TLXbar_io_in_0_a_bits_opcode;
  wire [2:0] TLXbar_io_in_0_a_bits_param;
  wire [3:0] TLXbar_io_in_0_a_bits_size;
  wire  TLXbar_io_in_0_a_bits_source;
  wire [31:0] TLXbar_io_in_0_a_bits_address;
  wire [3:0] TLXbar_io_in_0_a_bits_mask;
  wire [31:0] TLXbar_io_in_0_a_bits_data;
  wire  TLXbar_io_in_0_d_ready;
  wire  TLXbar_io_in_0_d_valid;
  wire [2:0] TLXbar_io_in_0_d_bits_opcode;
  wire [3:0] TLXbar_io_in_0_d_bits_size;
  wire  TLXbar_io_in_0_d_bits_source;
  wire [31:0] TLXbar_io_in_0_d_bits_data;
  wire  TLXbar_io_in_0_d_bits_error;
  wire  TLXbar_io_out_2_a_ready;
  wire  TLXbar_io_out_2_a_valid;
  wire [2:0] TLXbar_io_out_2_a_bits_opcode;
  wire [3:0] TLXbar_io_out_2_a_bits_size;
  wire [4:0] TLXbar_io_out_2_a_bits_source;
  wire  TLXbar_io_out_2_d_ready;
  wire  TLXbar_io_out_2_d_valid;
  wire [2:0] TLXbar_io_out_2_d_bits_opcode;
  wire [1:0] TLXbar_io_out_2_d_bits_param;
  wire [3:0] TLXbar_io_out_2_d_bits_size;
  wire [4:0] TLXbar_io_out_2_d_bits_source;
  wire  TLXbar_io_out_2_d_bits_sink;
  wire [31:0] TLXbar_io_out_2_d_bits_data;
  wire  TLXbar_io_out_2_d_bits_error;
  wire  TLXbar_io_out_1_a_ready;
  wire  TLXbar_io_out_1_a_valid;
  wire [2:0] TLXbar_io_out_1_a_bits_opcode;
  wire [3:0] TLXbar_io_out_1_a_bits_size;
  wire [4:0] TLXbar_io_out_1_a_bits_source;
  wire [30:0] TLXbar_io_out_1_a_bits_address;
  wire [3:0] TLXbar_io_out_1_a_bits_mask;
  wire [31:0] TLXbar_io_out_1_a_bits_data;
  wire  TLXbar_io_out_1_d_ready;
  wire  TLXbar_io_out_1_d_valid;
  wire [2:0] TLXbar_io_out_1_d_bits_opcode;
  wire [1:0] TLXbar_io_out_1_d_bits_param;
  wire [3:0] TLXbar_io_out_1_d_bits_size;
  wire [4:0] TLXbar_io_out_1_d_bits_source;
  wire  TLXbar_io_out_1_d_bits_sink;
  wire [31:0] TLXbar_io_out_1_d_bits_data;
  wire  TLXbar_io_out_1_d_bits_error;
  wire  TLXbar_io_out_0_a_ready;
  wire  TLXbar_io_out_0_a_valid;
  wire [2:0] TLXbar_io_out_0_a_bits_opcode;
  wire [2:0] TLXbar_io_out_0_a_bits_param;
  wire [2:0] TLXbar_io_out_0_a_bits_size;
  wire [4:0] TLXbar_io_out_0_a_bits_source;
  wire [31:0] TLXbar_io_out_0_a_bits_address;
  wire [3:0] TLXbar_io_out_0_a_bits_mask;
  wire [31:0] TLXbar_io_out_0_a_bits_data;
  wire  TLXbar_io_out_0_d_ready;
  wire  TLXbar_io_out_0_d_valid;
  wire [2:0] TLXbar_io_out_0_d_bits_opcode;
  wire [1:0] TLXbar_io_out_0_d_bits_param;
  wire [2:0] TLXbar_io_out_0_d_bits_size;
  wire [4:0] TLXbar_io_out_0_d_bits_source;
  wire  TLXbar_io_out_0_d_bits_sink;
  wire [31:0] TLXbar_io_out_0_d_bits_data;
  wire  TLXbar_io_out_0_d_bits_error;
  wire  TLBuffer_1_clock;
  wire  TLBuffer_1_reset;
  wire  TLBuffer_1_io_in_2_a_ready;
  wire  TLBuffer_1_io_in_2_a_valid;
  wire [2:0] TLBuffer_1_io_in_2_a_bits_opcode;
  wire [3:0] TLBuffer_1_io_in_2_a_bits_size;
  wire [4:0] TLBuffer_1_io_in_2_a_bits_source;
  wire  TLBuffer_1_io_in_2_d_ready;
  wire  TLBuffer_1_io_in_2_d_valid;
  wire [2:0] TLBuffer_1_io_in_2_d_bits_opcode;
  wire [1:0] TLBuffer_1_io_in_2_d_bits_param;
  wire [3:0] TLBuffer_1_io_in_2_d_bits_size;
  wire [4:0] TLBuffer_1_io_in_2_d_bits_source;
  wire  TLBuffer_1_io_in_2_d_bits_sink;
  wire [31:0] TLBuffer_1_io_in_2_d_bits_data;
  wire  TLBuffer_1_io_in_2_d_bits_error;
  wire  TLBuffer_1_io_in_1_a_ready;
  wire  TLBuffer_1_io_in_1_a_valid;
  wire [2:0] TLBuffer_1_io_in_1_a_bits_opcode;
  wire [3:0] TLBuffer_1_io_in_1_a_bits_size;
  wire [4:0] TLBuffer_1_io_in_1_a_bits_source;
  wire [30:0] TLBuffer_1_io_in_1_a_bits_address;
  wire [3:0] TLBuffer_1_io_in_1_a_bits_mask;
  wire [31:0] TLBuffer_1_io_in_1_a_bits_data;
  wire  TLBuffer_1_io_in_1_d_ready;
  wire  TLBuffer_1_io_in_1_d_valid;
  wire [2:0] TLBuffer_1_io_in_1_d_bits_opcode;
  wire [1:0] TLBuffer_1_io_in_1_d_bits_param;
  wire [3:0] TLBuffer_1_io_in_1_d_bits_size;
  wire [4:0] TLBuffer_1_io_in_1_d_bits_source;
  wire  TLBuffer_1_io_in_1_d_bits_sink;
  wire [31:0] TLBuffer_1_io_in_1_d_bits_data;
  wire  TLBuffer_1_io_in_1_d_bits_error;
  wire  TLBuffer_1_io_in_0_a_ready;
  wire  TLBuffer_1_io_in_0_a_valid;
  wire [2:0] TLBuffer_1_io_in_0_a_bits_opcode;
  wire [2:0] TLBuffer_1_io_in_0_a_bits_param;
  wire [2:0] TLBuffer_1_io_in_0_a_bits_size;
  wire [4:0] TLBuffer_1_io_in_0_a_bits_source;
  wire [31:0] TLBuffer_1_io_in_0_a_bits_address;
  wire [3:0] TLBuffer_1_io_in_0_a_bits_mask;
  wire [31:0] TLBuffer_1_io_in_0_a_bits_data;
  wire  TLBuffer_1_io_in_0_d_ready;
  wire  TLBuffer_1_io_in_0_d_valid;
  wire [2:0] TLBuffer_1_io_in_0_d_bits_opcode;
  wire [1:0] TLBuffer_1_io_in_0_d_bits_param;
  wire [2:0] TLBuffer_1_io_in_0_d_bits_size;
  wire [4:0] TLBuffer_1_io_in_0_d_bits_source;
  wire  TLBuffer_1_io_in_0_d_bits_sink;
  wire [31:0] TLBuffer_1_io_in_0_d_bits_data;
  wire  TLBuffer_1_io_in_0_d_bits_error;
  wire  TLBuffer_1_io_out_2_a_ready;
  wire  TLBuffer_1_io_out_2_a_valid;
  wire [2:0] TLBuffer_1_io_out_2_a_bits_opcode;
  wire [3:0] TLBuffer_1_io_out_2_a_bits_size;
  wire [4:0] TLBuffer_1_io_out_2_a_bits_source;
  wire  TLBuffer_1_io_out_2_d_ready;
  wire  TLBuffer_1_io_out_2_d_valid;
  wire [2:0] TLBuffer_1_io_out_2_d_bits_opcode;
  wire [1:0] TLBuffer_1_io_out_2_d_bits_param;
  wire [3:0] TLBuffer_1_io_out_2_d_bits_size;
  wire [4:0] TLBuffer_1_io_out_2_d_bits_source;
  wire  TLBuffer_1_io_out_2_d_bits_sink;
  wire [31:0] TLBuffer_1_io_out_2_d_bits_data;
  wire  TLBuffer_1_io_out_2_d_bits_error;
  wire  TLBuffer_1_io_out_1_a_ready;
  wire  TLBuffer_1_io_out_1_a_valid;
  wire [2:0] TLBuffer_1_io_out_1_a_bits_opcode;
  wire [3:0] TLBuffer_1_io_out_1_a_bits_size;
  wire [4:0] TLBuffer_1_io_out_1_a_bits_source;
  wire [30:0] TLBuffer_1_io_out_1_a_bits_address;
  wire [3:0] TLBuffer_1_io_out_1_a_bits_mask;
  wire [31:0] TLBuffer_1_io_out_1_a_bits_data;
  wire  TLBuffer_1_io_out_1_d_ready;
  wire  TLBuffer_1_io_out_1_d_valid;
  wire [2:0] TLBuffer_1_io_out_1_d_bits_opcode;
  wire [1:0] TLBuffer_1_io_out_1_d_bits_param;
  wire [3:0] TLBuffer_1_io_out_1_d_bits_size;
  wire [4:0] TLBuffer_1_io_out_1_d_bits_source;
  wire  TLBuffer_1_io_out_1_d_bits_sink;
  wire [31:0] TLBuffer_1_io_out_1_d_bits_data;
  wire  TLBuffer_1_io_out_1_d_bits_error;
  wire  TLBuffer_1_io_out_0_a_ready;
  wire  TLBuffer_1_io_out_0_a_valid;
  wire [2:0] TLBuffer_1_io_out_0_a_bits_opcode;
  wire [2:0] TLBuffer_1_io_out_0_a_bits_param;
  wire [2:0] TLBuffer_1_io_out_0_a_bits_size;
  wire [4:0] TLBuffer_1_io_out_0_a_bits_source;
  wire [31:0] TLBuffer_1_io_out_0_a_bits_address;
  wire [3:0] TLBuffer_1_io_out_0_a_bits_mask;
  wire [31:0] TLBuffer_1_io_out_0_a_bits_data;
  wire  TLBuffer_1_io_out_0_d_ready;
  wire  TLBuffer_1_io_out_0_d_valid;
  wire [2:0] TLBuffer_1_io_out_0_d_bits_opcode;
  wire [1:0] TLBuffer_1_io_out_0_d_bits_param;
  wire [2:0] TLBuffer_1_io_out_0_d_bits_size;
  wire [4:0] TLBuffer_1_io_out_0_d_bits_source;
  wire  TLBuffer_1_io_out_0_d_bits_sink;
  wire [31:0] TLBuffer_1_io_out_0_d_bits_data;
  wire  TLBuffer_1_io_out_0_d_bits_error;
  wire  TLWidthWidget_clock;
  wire  TLWidthWidget_reset;
  wire  TLWidthWidget_io_in_1_a_ready;
  wire  TLWidthWidget_io_in_1_a_valid;
  wire [2:0] TLWidthWidget_io_in_1_a_bits_opcode;
  wire [3:0] TLWidthWidget_io_in_1_a_bits_size;
  wire [4:0] TLWidthWidget_io_in_1_a_bits_source;
  wire [30:0] TLWidthWidget_io_in_1_a_bits_address;
  wire [3:0] TLWidthWidget_io_in_1_a_bits_mask;
  wire [31:0] TLWidthWidget_io_in_1_a_bits_data;
  wire  TLWidthWidget_io_in_1_d_ready;
  wire  TLWidthWidget_io_in_1_d_valid;
  wire [2:0] TLWidthWidget_io_in_1_d_bits_opcode;
  wire [1:0] TLWidthWidget_io_in_1_d_bits_param;
  wire [3:0] TLWidthWidget_io_in_1_d_bits_size;
  wire [4:0] TLWidthWidget_io_in_1_d_bits_source;
  wire  TLWidthWidget_io_in_1_d_bits_sink;
  wire [31:0] TLWidthWidget_io_in_1_d_bits_data;
  wire  TLWidthWidget_io_in_1_d_bits_error;
  wire  TLWidthWidget_io_in_0_a_ready;
  wire  TLWidthWidget_io_in_0_a_valid;
  wire [2:0] TLWidthWidget_io_in_0_a_bits_opcode;
  wire [2:0] TLWidthWidget_io_in_0_a_bits_param;
  wire [2:0] TLWidthWidget_io_in_0_a_bits_size;
  wire [4:0] TLWidthWidget_io_in_0_a_bits_source;
  wire [31:0] TLWidthWidget_io_in_0_a_bits_address;
  wire [3:0] TLWidthWidget_io_in_0_a_bits_mask;
  wire [31:0] TLWidthWidget_io_in_0_a_bits_data;
  wire  TLWidthWidget_io_in_0_d_ready;
  wire  TLWidthWidget_io_in_0_d_valid;
  wire [2:0] TLWidthWidget_io_in_0_d_bits_opcode;
  wire [1:0] TLWidthWidget_io_in_0_d_bits_param;
  wire [2:0] TLWidthWidget_io_in_0_d_bits_size;
  wire [4:0] TLWidthWidget_io_in_0_d_bits_source;
  wire  TLWidthWidget_io_in_0_d_bits_sink;
  wire [31:0] TLWidthWidget_io_in_0_d_bits_data;
  wire  TLWidthWidget_io_in_0_d_bits_error;
  wire  TLWidthWidget_io_out_1_a_ready;
  wire  TLWidthWidget_io_out_1_a_valid;
  wire [2:0] TLWidthWidget_io_out_1_a_bits_opcode;
  wire [3:0] TLWidthWidget_io_out_1_a_bits_size;
  wire [4:0] TLWidthWidget_io_out_1_a_bits_source;
  wire [30:0] TLWidthWidget_io_out_1_a_bits_address;
  wire [7:0] TLWidthWidget_io_out_1_a_bits_mask;
  wire [63:0] TLWidthWidget_io_out_1_a_bits_data;
  wire  TLWidthWidget_io_out_1_d_ready;
  wire  TLWidthWidget_io_out_1_d_valid;
  wire [2:0] TLWidthWidget_io_out_1_d_bits_opcode;
  wire [1:0] TLWidthWidget_io_out_1_d_bits_param;
  wire [3:0] TLWidthWidget_io_out_1_d_bits_size;
  wire [4:0] TLWidthWidget_io_out_1_d_bits_source;
  wire  TLWidthWidget_io_out_1_d_bits_sink;
  wire [63:0] TLWidthWidget_io_out_1_d_bits_data;
  wire  TLWidthWidget_io_out_1_d_bits_error;
  wire  TLWidthWidget_io_out_0_a_ready;
  wire  TLWidthWidget_io_out_0_a_valid;
  wire [2:0] TLWidthWidget_io_out_0_a_bits_opcode;
  wire [2:0] TLWidthWidget_io_out_0_a_bits_param;
  wire [2:0] TLWidthWidget_io_out_0_a_bits_size;
  wire [4:0] TLWidthWidget_io_out_0_a_bits_source;
  wire [31:0] TLWidthWidget_io_out_0_a_bits_address;
  wire [3:0] TLWidthWidget_io_out_0_a_bits_mask;
  wire [31:0] TLWidthWidget_io_out_0_a_bits_data;
  wire  TLWidthWidget_io_out_0_d_ready;
  wire  TLWidthWidget_io_out_0_d_valid;
  wire [2:0] TLWidthWidget_io_out_0_d_bits_opcode;
  wire [1:0] TLWidthWidget_io_out_0_d_bits_param;
  wire [2:0] TLWidthWidget_io_out_0_d_bits_size;
  wire [4:0] TLWidthWidget_io_out_0_d_bits_source;
  wire  TLWidthWidget_io_out_0_d_bits_sink;
  wire [31:0] TLWidthWidget_io_out_0_d_bits_data;
  wire  TLWidthWidget_io_out_0_d_bits_error;
  wire  TLSplitter_io_in_1_a_ready;
  wire  TLSplitter_io_in_1_a_valid;
  wire [2:0] TLSplitter_io_in_1_a_bits_opcode;
  wire [2:0] TLSplitter_io_in_1_a_bits_param;
  wire [3:0] TLSplitter_io_in_1_a_bits_size;
  wire [3:0] TLSplitter_io_in_1_a_bits_source;
  wire [31:0] TLSplitter_io_in_1_a_bits_address;
  wire [3:0] TLSplitter_io_in_1_a_bits_mask;
  wire [31:0] TLSplitter_io_in_1_a_bits_data;
  wire  TLSplitter_io_in_1_d_ready;
  wire  TLSplitter_io_in_1_d_valid;
  wire [2:0] TLSplitter_io_in_1_d_bits_opcode;
  wire [3:0] TLSplitter_io_in_1_d_bits_size;
  wire [3:0] TLSplitter_io_in_1_d_bits_source;
  wire  TLSplitter_io_in_0_a_ready;
  wire  TLSplitter_io_in_0_a_valid;
  wire [2:0] TLSplitter_io_in_0_a_bits_opcode;
  wire [2:0] TLSplitter_io_in_0_a_bits_param;
  wire [3:0] TLSplitter_io_in_0_a_bits_size;
  wire  TLSplitter_io_in_0_a_bits_source;
  wire [31:0] TLSplitter_io_in_0_a_bits_address;
  wire [3:0] TLSplitter_io_in_0_a_bits_mask;
  wire [31:0] TLSplitter_io_in_0_a_bits_data;
  wire  TLSplitter_io_in_0_d_ready;
  wire  TLSplitter_io_in_0_d_valid;
  wire [2:0] TLSplitter_io_in_0_d_bits_opcode;
  wire [3:0] TLSplitter_io_in_0_d_bits_size;
  wire  TLSplitter_io_in_0_d_bits_source;
  wire [31:0] TLSplitter_io_in_0_d_bits_data;
  wire  TLSplitter_io_in_0_d_bits_error;
  wire  TLSplitter_io_out_1_a_ready;
  wire  TLSplitter_io_out_1_a_valid;
  wire [2:0] TLSplitter_io_out_1_a_bits_opcode;
  wire [2:0] TLSplitter_io_out_1_a_bits_param;
  wire [3:0] TLSplitter_io_out_1_a_bits_size;
  wire [3:0] TLSplitter_io_out_1_a_bits_source;
  wire [31:0] TLSplitter_io_out_1_a_bits_address;
  wire [3:0] TLSplitter_io_out_1_a_bits_mask;
  wire [31:0] TLSplitter_io_out_1_a_bits_data;
  wire  TLSplitter_io_out_1_d_ready;
  wire  TLSplitter_io_out_1_d_valid;
  wire [2:0] TLSplitter_io_out_1_d_bits_opcode;
  wire [3:0] TLSplitter_io_out_1_d_bits_size;
  wire [3:0] TLSplitter_io_out_1_d_bits_source;
  wire  TLSplitter_io_out_0_a_ready;
  wire  TLSplitter_io_out_0_a_valid;
  wire [2:0] TLSplitter_io_out_0_a_bits_opcode;
  wire [2:0] TLSplitter_io_out_0_a_bits_param;
  wire [3:0] TLSplitter_io_out_0_a_bits_size;
  wire  TLSplitter_io_out_0_a_bits_source;
  wire [31:0] TLSplitter_io_out_0_a_bits_address;
  wire [3:0] TLSplitter_io_out_0_a_bits_mask;
  wire [31:0] TLSplitter_io_out_0_a_bits_data;
  wire  TLSplitter_io_out_0_d_ready;
  wire  TLSplitter_io_out_0_d_valid;
  wire [2:0] TLSplitter_io_out_0_d_bits_opcode;
  wire [3:0] TLSplitter_io_out_0_d_bits_size;
  wire  TLSplitter_io_out_0_d_bits_source;
  wire [31:0] TLSplitter_io_out_0_d_bits_data;
  wire  TLSplitter_io_out_0_d_bits_error;
  wire  TLFIFOFixer_io_in_0_a_ready;
  wire  TLFIFOFixer_io_in_0_a_valid;
  wire [2:0] TLFIFOFixer_io_in_0_a_bits_opcode;
  wire [2:0] TLFIFOFixer_io_in_0_a_bits_param;
  wire [3:0] TLFIFOFixer_io_in_0_a_bits_size;
  wire  TLFIFOFixer_io_in_0_a_bits_source;
  wire [31:0] TLFIFOFixer_io_in_0_a_bits_address;
  wire [3:0] TLFIFOFixer_io_in_0_a_bits_mask;
  wire [31:0] TLFIFOFixer_io_in_0_a_bits_data;
  wire  TLFIFOFixer_io_in_0_d_ready;
  wire  TLFIFOFixer_io_in_0_d_valid;
  wire [2:0] TLFIFOFixer_io_in_0_d_bits_opcode;
  wire [3:0] TLFIFOFixer_io_in_0_d_bits_size;
  wire  TLFIFOFixer_io_in_0_d_bits_source;
  wire [31:0] TLFIFOFixer_io_in_0_d_bits_data;
  wire  TLFIFOFixer_io_in_0_d_bits_error;
  wire  TLFIFOFixer_io_out_0_a_ready;
  wire  TLFIFOFixer_io_out_0_a_valid;
  wire [2:0] TLFIFOFixer_io_out_0_a_bits_opcode;
  wire [2:0] TLFIFOFixer_io_out_0_a_bits_param;
  wire [3:0] TLFIFOFixer_io_out_0_a_bits_size;
  wire  TLFIFOFixer_io_out_0_a_bits_source;
  wire [31:0] TLFIFOFixer_io_out_0_a_bits_address;
  wire [3:0] TLFIFOFixer_io_out_0_a_bits_mask;
  wire [31:0] TLFIFOFixer_io_out_0_a_bits_data;
  wire  TLFIFOFixer_io_out_0_d_ready;
  wire  TLFIFOFixer_io_out_0_d_valid;
  wire [2:0] TLFIFOFixer_io_out_0_d_bits_opcode;
  wire [3:0] TLFIFOFixer_io_out_0_d_bits_size;
  wire  TLFIFOFixer_io_out_0_d_bits_source;
  wire [31:0] TLFIFOFixer_io_out_0_d_bits_data;
  wire  TLFIFOFixer_io_out_0_d_bits_error;
  wire  TLFIFOFixer_1_clock;
  wire  TLFIFOFixer_1_reset;
  wire  TLFIFOFixer_1_io_in_0_a_ready;
  wire  TLFIFOFixer_1_io_in_0_a_valid;
  wire [2:0] TLFIFOFixer_1_io_in_0_a_bits_opcode;
  wire [2:0] TLFIFOFixer_1_io_in_0_a_bits_param;
  wire [3:0] TLFIFOFixer_1_io_in_0_a_bits_size;
  wire [3:0] TLFIFOFixer_1_io_in_0_a_bits_source;
  wire [31:0] TLFIFOFixer_1_io_in_0_a_bits_address;
  wire [3:0] TLFIFOFixer_1_io_in_0_a_bits_mask;
  wire [31:0] TLFIFOFixer_1_io_in_0_a_bits_data;
  wire  TLFIFOFixer_1_io_in_0_d_ready;
  wire  TLFIFOFixer_1_io_in_0_d_valid;
  wire [2:0] TLFIFOFixer_1_io_in_0_d_bits_opcode;
  wire [3:0] TLFIFOFixer_1_io_in_0_d_bits_size;
  wire [3:0] TLFIFOFixer_1_io_in_0_d_bits_source;
  wire  TLFIFOFixer_1_io_out_0_a_ready;
  wire  TLFIFOFixer_1_io_out_0_a_valid;
  wire [2:0] TLFIFOFixer_1_io_out_0_a_bits_opcode;
  wire [2:0] TLFIFOFixer_1_io_out_0_a_bits_param;
  wire [3:0] TLFIFOFixer_1_io_out_0_a_bits_size;
  wire [3:0] TLFIFOFixer_1_io_out_0_a_bits_source;
  wire [31:0] TLFIFOFixer_1_io_out_0_a_bits_address;
  wire [3:0] TLFIFOFixer_1_io_out_0_a_bits_mask;
  wire [31:0] TLFIFOFixer_1_io_out_0_a_bits_data;
  wire  TLFIFOFixer_1_io_out_0_d_ready;
  wire  TLFIFOFixer_1_io_out_0_d_valid;
  wire [2:0] TLFIFOFixer_1_io_out_0_d_bits_opcode;
  wire [3:0] TLFIFOFixer_1_io_out_0_d_bits_size;
  wire [3:0] TLFIFOFixer_1_io_out_0_d_bits_source;
  wire  TLXbar_1_clock;
  wire  TLXbar_1_reset;
  wire  TLXbar_1_io_in_0_a_ready;
  wire  TLXbar_1_io_in_0_a_valid;
  wire [2:0] TLXbar_1_io_in_0_a_bits_opcode;
  wire [2:0] TLXbar_1_io_in_0_a_bits_param;
  wire [2:0] TLXbar_1_io_in_0_a_bits_size;
  wire [4:0] TLXbar_1_io_in_0_a_bits_source;
  wire [31:0] TLXbar_1_io_in_0_a_bits_address;
  wire [3:0] TLXbar_1_io_in_0_a_bits_mask;
  wire [31:0] TLXbar_1_io_in_0_a_bits_data;
  wire  TLXbar_1_io_in_0_d_ready;
  wire  TLXbar_1_io_in_0_d_valid;
  wire [2:0] TLXbar_1_io_in_0_d_bits_opcode;
  wire [1:0] TLXbar_1_io_in_0_d_bits_param;
  wire [2:0] TLXbar_1_io_in_0_d_bits_size;
  wire [4:0] TLXbar_1_io_in_0_d_bits_source;
  wire  TLXbar_1_io_in_0_d_bits_sink;
  wire [31:0] TLXbar_1_io_in_0_d_bits_data;
  wire  TLXbar_1_io_in_0_d_bits_error;
  wire  TLXbar_1_io_out_4_a_ready;
  wire  TLXbar_1_io_out_4_a_valid;
  wire [2:0] TLXbar_1_io_out_4_a_bits_opcode;
  wire [2:0] TLXbar_1_io_out_4_a_bits_param;
  wire [2:0] TLXbar_1_io_out_4_a_bits_size;
  wire [4:0] TLXbar_1_io_out_4_a_bits_source;
  wire [31:0] TLXbar_1_io_out_4_a_bits_address;
  wire [3:0] TLXbar_1_io_out_4_a_bits_mask;
  wire [31:0] TLXbar_1_io_out_4_a_bits_data;
  wire  TLXbar_1_io_out_4_d_ready;
  wire  TLXbar_1_io_out_4_d_valid;
  wire [2:0] TLXbar_1_io_out_4_d_bits_opcode;
  wire [1:0] TLXbar_1_io_out_4_d_bits_param;
  wire [2:0] TLXbar_1_io_out_4_d_bits_size;
  wire [4:0] TLXbar_1_io_out_4_d_bits_source;
  wire  TLXbar_1_io_out_4_d_bits_sink;
  wire [31:0] TLXbar_1_io_out_4_d_bits_data;
  wire  TLXbar_1_io_out_4_d_bits_error;
  wire  TLXbar_1_io_out_3_a_ready;
  wire  TLXbar_1_io_out_3_a_valid;
  wire [2:0] TLXbar_1_io_out_3_a_bits_opcode;
  wire [2:0] TLXbar_1_io_out_3_a_bits_size;
  wire [4:0] TLXbar_1_io_out_3_a_bits_source;
  wire [16:0] TLXbar_1_io_out_3_a_bits_address;
  wire [3:0] TLXbar_1_io_out_3_a_bits_mask;
  wire  TLXbar_1_io_out_3_d_ready;
  wire  TLXbar_1_io_out_3_d_valid;
  wire [2:0] TLXbar_1_io_out_3_d_bits_opcode;
  wire [1:0] TLXbar_1_io_out_3_d_bits_param;
  wire [2:0] TLXbar_1_io_out_3_d_bits_size;
  wire [4:0] TLXbar_1_io_out_3_d_bits_source;
  wire  TLXbar_1_io_out_3_d_bits_sink;
  wire [31:0] TLXbar_1_io_out_3_d_bits_data;
  wire  TLXbar_1_io_out_3_d_bits_error;
  wire  TLXbar_1_io_out_2_a_ready;
  wire  TLXbar_1_io_out_2_a_valid;
  wire [2:0] TLXbar_1_io_out_2_a_bits_opcode;
  wire [2:0] TLXbar_1_io_out_2_a_bits_size;
  wire [4:0] TLXbar_1_io_out_2_a_bits_source;
  wire [11:0] TLXbar_1_io_out_2_a_bits_address;
  wire [3:0] TLXbar_1_io_out_2_a_bits_mask;
  wire [31:0] TLXbar_1_io_out_2_a_bits_data;
  wire  TLXbar_1_io_out_2_d_ready;
  wire  TLXbar_1_io_out_2_d_valid;
  wire [2:0] TLXbar_1_io_out_2_d_bits_opcode;
  wire [1:0] TLXbar_1_io_out_2_d_bits_param;
  wire [2:0] TLXbar_1_io_out_2_d_bits_size;
  wire [4:0] TLXbar_1_io_out_2_d_bits_source;
  wire  TLXbar_1_io_out_2_d_bits_sink;
  wire [31:0] TLXbar_1_io_out_2_d_bits_data;
  wire  TLXbar_1_io_out_2_d_bits_error;
  wire  TLXbar_1_io_out_1_a_ready;
  wire  TLXbar_1_io_out_1_a_valid;
  wire [2:0] TLXbar_1_io_out_1_a_bits_opcode;
  wire [2:0] TLXbar_1_io_out_1_a_bits_size;
  wire [4:0] TLXbar_1_io_out_1_a_bits_source;
  wire [25:0] TLXbar_1_io_out_1_a_bits_address;
  wire [3:0] TLXbar_1_io_out_1_a_bits_mask;
  wire [31:0] TLXbar_1_io_out_1_a_bits_data;
  wire  TLXbar_1_io_out_1_d_ready;
  wire  TLXbar_1_io_out_1_d_valid;
  wire [2:0] TLXbar_1_io_out_1_d_bits_opcode;
  wire [1:0] TLXbar_1_io_out_1_d_bits_param;
  wire [2:0] TLXbar_1_io_out_1_d_bits_size;
  wire [4:0] TLXbar_1_io_out_1_d_bits_source;
  wire  TLXbar_1_io_out_1_d_bits_sink;
  wire [31:0] TLXbar_1_io_out_1_d_bits_data;
  wire  TLXbar_1_io_out_1_d_bits_error;
  wire  TLXbar_1_io_out_0_a_ready;
  wire  TLXbar_1_io_out_0_a_valid;
  wire [2:0] TLXbar_1_io_out_0_a_bits_opcode;
  wire [2:0] TLXbar_1_io_out_0_a_bits_size;
  wire [4:0] TLXbar_1_io_out_0_a_bits_source;
  wire [27:0] TLXbar_1_io_out_0_a_bits_address;
  wire [3:0] TLXbar_1_io_out_0_a_bits_mask;
  wire [31:0] TLXbar_1_io_out_0_a_bits_data;
  wire  TLXbar_1_io_out_0_d_ready;
  wire  TLXbar_1_io_out_0_d_valid;
  wire [2:0] TLXbar_1_io_out_0_d_bits_opcode;
  wire [1:0] TLXbar_1_io_out_0_d_bits_param;
  wire [2:0] TLXbar_1_io_out_0_d_bits_size;
  wire [4:0] TLXbar_1_io_out_0_d_bits_source;
  wire  TLXbar_1_io_out_0_d_bits_sink;
  wire [31:0] TLXbar_1_io_out_0_d_bits_data;
  wire  TLXbar_1_io_out_0_d_bits_error;
  wire  TLBuffer_2_clock;
  wire  TLBuffer_2_reset;
  wire  TLBuffer_2_io_in_0_a_ready;
  wire  TLBuffer_2_io_in_0_a_valid;
  wire [2:0] TLBuffer_2_io_in_0_a_bits_opcode;
  wire [2:0] TLBuffer_2_io_in_0_a_bits_param;
  wire [2:0] TLBuffer_2_io_in_0_a_bits_size;
  wire [4:0] TLBuffer_2_io_in_0_a_bits_source;
  wire [31:0] TLBuffer_2_io_in_0_a_bits_address;
  wire [3:0] TLBuffer_2_io_in_0_a_bits_mask;
  wire [31:0] TLBuffer_2_io_in_0_a_bits_data;
  wire  TLBuffer_2_io_in_0_d_ready;
  wire  TLBuffer_2_io_in_0_d_valid;
  wire [2:0] TLBuffer_2_io_in_0_d_bits_opcode;
  wire [1:0] TLBuffer_2_io_in_0_d_bits_param;
  wire [2:0] TLBuffer_2_io_in_0_d_bits_size;
  wire [4:0] TLBuffer_2_io_in_0_d_bits_source;
  wire  TLBuffer_2_io_in_0_d_bits_sink;
  wire [31:0] TLBuffer_2_io_in_0_d_bits_data;
  wire  TLBuffer_2_io_in_0_d_bits_error;
  wire  TLBuffer_2_io_out_0_a_ready;
  wire  TLBuffer_2_io_out_0_a_valid;
  wire [2:0] TLBuffer_2_io_out_0_a_bits_opcode;
  wire [2:0] TLBuffer_2_io_out_0_a_bits_param;
  wire [2:0] TLBuffer_2_io_out_0_a_bits_size;
  wire [4:0] TLBuffer_2_io_out_0_a_bits_source;
  wire [31:0] TLBuffer_2_io_out_0_a_bits_address;
  wire [3:0] TLBuffer_2_io_out_0_a_bits_mask;
  wire [31:0] TLBuffer_2_io_out_0_a_bits_data;
  wire  TLBuffer_2_io_out_0_d_ready;
  wire  TLBuffer_2_io_out_0_d_valid;
  wire [2:0] TLBuffer_2_io_out_0_d_bits_opcode;
  wire [1:0] TLBuffer_2_io_out_0_d_bits_param;
  wire [2:0] TLBuffer_2_io_out_0_d_bits_size;
  wire [4:0] TLBuffer_2_io_out_0_d_bits_source;
  wire  TLBuffer_2_io_out_0_d_bits_sink;
  wire [31:0] TLBuffer_2_io_out_0_d_bits_data;
  wire  TLBuffer_2_io_out_0_d_bits_error;
  wire  TLBuffer_3_io_in_4_a_ready;
  wire  TLBuffer_3_io_in_4_a_valid;
  wire [2:0] TLBuffer_3_io_in_4_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_in_4_a_bits_param;
  wire [2:0] TLBuffer_3_io_in_4_a_bits_size;
  wire [4:0] TLBuffer_3_io_in_4_a_bits_source;
  wire [31:0] TLBuffer_3_io_in_4_a_bits_address;
  wire [3:0] TLBuffer_3_io_in_4_a_bits_mask;
  wire [31:0] TLBuffer_3_io_in_4_a_bits_data;
  wire  TLBuffer_3_io_in_4_d_ready;
  wire  TLBuffer_3_io_in_4_d_valid;
  wire [2:0] TLBuffer_3_io_in_4_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_in_4_d_bits_param;
  wire [2:0] TLBuffer_3_io_in_4_d_bits_size;
  wire [4:0] TLBuffer_3_io_in_4_d_bits_source;
  wire  TLBuffer_3_io_in_4_d_bits_sink;
  wire [31:0] TLBuffer_3_io_in_4_d_bits_data;
  wire  TLBuffer_3_io_in_4_d_bits_error;
  wire  TLBuffer_3_io_in_3_a_ready;
  wire  TLBuffer_3_io_in_3_a_valid;
  wire [2:0] TLBuffer_3_io_in_3_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_in_3_a_bits_size;
  wire [4:0] TLBuffer_3_io_in_3_a_bits_source;
  wire [16:0] TLBuffer_3_io_in_3_a_bits_address;
  wire [3:0] TLBuffer_3_io_in_3_a_bits_mask;
  wire  TLBuffer_3_io_in_3_d_ready;
  wire  TLBuffer_3_io_in_3_d_valid;
  wire [2:0] TLBuffer_3_io_in_3_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_in_3_d_bits_param;
  wire [2:0] TLBuffer_3_io_in_3_d_bits_size;
  wire [4:0] TLBuffer_3_io_in_3_d_bits_source;
  wire  TLBuffer_3_io_in_3_d_bits_sink;
  wire [31:0] TLBuffer_3_io_in_3_d_bits_data;
  wire  TLBuffer_3_io_in_3_d_bits_error;
  wire  TLBuffer_3_io_in_2_a_ready;
  wire  TLBuffer_3_io_in_2_a_valid;
  wire [2:0] TLBuffer_3_io_in_2_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_in_2_a_bits_size;
  wire [4:0] TLBuffer_3_io_in_2_a_bits_source;
  wire [11:0] TLBuffer_3_io_in_2_a_bits_address;
  wire [3:0] TLBuffer_3_io_in_2_a_bits_mask;
  wire [31:0] TLBuffer_3_io_in_2_a_bits_data;
  wire  TLBuffer_3_io_in_2_d_ready;
  wire  TLBuffer_3_io_in_2_d_valid;
  wire [2:0] TLBuffer_3_io_in_2_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_in_2_d_bits_param;
  wire [2:0] TLBuffer_3_io_in_2_d_bits_size;
  wire [4:0] TLBuffer_3_io_in_2_d_bits_source;
  wire  TLBuffer_3_io_in_2_d_bits_sink;
  wire [31:0] TLBuffer_3_io_in_2_d_bits_data;
  wire  TLBuffer_3_io_in_2_d_bits_error;
  wire  TLBuffer_3_io_in_1_a_ready;
  wire  TLBuffer_3_io_in_1_a_valid;
  wire [2:0] TLBuffer_3_io_in_1_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_in_1_a_bits_size;
  wire [4:0] TLBuffer_3_io_in_1_a_bits_source;
  wire [25:0] TLBuffer_3_io_in_1_a_bits_address;
  wire [3:0] TLBuffer_3_io_in_1_a_bits_mask;
  wire [31:0] TLBuffer_3_io_in_1_a_bits_data;
  wire  TLBuffer_3_io_in_1_d_ready;
  wire  TLBuffer_3_io_in_1_d_valid;
  wire [2:0] TLBuffer_3_io_in_1_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_in_1_d_bits_param;
  wire [2:0] TLBuffer_3_io_in_1_d_bits_size;
  wire [4:0] TLBuffer_3_io_in_1_d_bits_source;
  wire  TLBuffer_3_io_in_1_d_bits_sink;
  wire [31:0] TLBuffer_3_io_in_1_d_bits_data;
  wire  TLBuffer_3_io_in_1_d_bits_error;
  wire  TLBuffer_3_io_in_0_a_ready;
  wire  TLBuffer_3_io_in_0_a_valid;
  wire [2:0] TLBuffer_3_io_in_0_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_in_0_a_bits_size;
  wire [4:0] TLBuffer_3_io_in_0_a_bits_source;
  wire [27:0] TLBuffer_3_io_in_0_a_bits_address;
  wire [3:0] TLBuffer_3_io_in_0_a_bits_mask;
  wire [31:0] TLBuffer_3_io_in_0_a_bits_data;
  wire  TLBuffer_3_io_in_0_d_ready;
  wire  TLBuffer_3_io_in_0_d_valid;
  wire [2:0] TLBuffer_3_io_in_0_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_in_0_d_bits_param;
  wire [2:0] TLBuffer_3_io_in_0_d_bits_size;
  wire [4:0] TLBuffer_3_io_in_0_d_bits_source;
  wire  TLBuffer_3_io_in_0_d_bits_sink;
  wire [31:0] TLBuffer_3_io_in_0_d_bits_data;
  wire  TLBuffer_3_io_in_0_d_bits_error;
  wire  TLBuffer_3_io_out_4_a_ready;
  wire  TLBuffer_3_io_out_4_a_valid;
  wire [2:0] TLBuffer_3_io_out_4_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_out_4_a_bits_param;
  wire [2:0] TLBuffer_3_io_out_4_a_bits_size;
  wire [4:0] TLBuffer_3_io_out_4_a_bits_source;
  wire [31:0] TLBuffer_3_io_out_4_a_bits_address;
  wire [3:0] TLBuffer_3_io_out_4_a_bits_mask;
  wire [31:0] TLBuffer_3_io_out_4_a_bits_data;
  wire  TLBuffer_3_io_out_4_d_ready;
  wire  TLBuffer_3_io_out_4_d_valid;
  wire [2:0] TLBuffer_3_io_out_4_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_out_4_d_bits_param;
  wire [2:0] TLBuffer_3_io_out_4_d_bits_size;
  wire [4:0] TLBuffer_3_io_out_4_d_bits_source;
  wire  TLBuffer_3_io_out_4_d_bits_sink;
  wire [31:0] TLBuffer_3_io_out_4_d_bits_data;
  wire  TLBuffer_3_io_out_4_d_bits_error;
  wire  TLBuffer_3_io_out_3_a_ready;
  wire  TLBuffer_3_io_out_3_a_valid;
  wire [2:0] TLBuffer_3_io_out_3_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_out_3_a_bits_size;
  wire [4:0] TLBuffer_3_io_out_3_a_bits_source;
  wire [16:0] TLBuffer_3_io_out_3_a_bits_address;
  wire [3:0] TLBuffer_3_io_out_3_a_bits_mask;
  wire  TLBuffer_3_io_out_3_d_ready;
  wire  TLBuffer_3_io_out_3_d_valid;
  wire [2:0] TLBuffer_3_io_out_3_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_out_3_d_bits_param;
  wire [2:0] TLBuffer_3_io_out_3_d_bits_size;
  wire [4:0] TLBuffer_3_io_out_3_d_bits_source;
  wire  TLBuffer_3_io_out_3_d_bits_sink;
  wire [31:0] TLBuffer_3_io_out_3_d_bits_data;
  wire  TLBuffer_3_io_out_3_d_bits_error;
  wire  TLBuffer_3_io_out_2_a_ready;
  wire  TLBuffer_3_io_out_2_a_valid;
  wire [2:0] TLBuffer_3_io_out_2_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_out_2_a_bits_size;
  wire [4:0] TLBuffer_3_io_out_2_a_bits_source;
  wire [11:0] TLBuffer_3_io_out_2_a_bits_address;
  wire [3:0] TLBuffer_3_io_out_2_a_bits_mask;
  wire [31:0] TLBuffer_3_io_out_2_a_bits_data;
  wire  TLBuffer_3_io_out_2_d_ready;
  wire  TLBuffer_3_io_out_2_d_valid;
  wire [2:0] TLBuffer_3_io_out_2_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_out_2_d_bits_param;
  wire [2:0] TLBuffer_3_io_out_2_d_bits_size;
  wire [4:0] TLBuffer_3_io_out_2_d_bits_source;
  wire  TLBuffer_3_io_out_2_d_bits_sink;
  wire [31:0] TLBuffer_3_io_out_2_d_bits_data;
  wire  TLBuffer_3_io_out_2_d_bits_error;
  wire  TLBuffer_3_io_out_1_a_ready;
  wire  TLBuffer_3_io_out_1_a_valid;
  wire [2:0] TLBuffer_3_io_out_1_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_out_1_a_bits_size;
  wire [4:0] TLBuffer_3_io_out_1_a_bits_source;
  wire [25:0] TLBuffer_3_io_out_1_a_bits_address;
  wire [3:0] TLBuffer_3_io_out_1_a_bits_mask;
  wire [31:0] TLBuffer_3_io_out_1_a_bits_data;
  wire  TLBuffer_3_io_out_1_d_ready;
  wire  TLBuffer_3_io_out_1_d_valid;
  wire [2:0] TLBuffer_3_io_out_1_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_out_1_d_bits_param;
  wire [2:0] TLBuffer_3_io_out_1_d_bits_size;
  wire [4:0] TLBuffer_3_io_out_1_d_bits_source;
  wire  TLBuffer_3_io_out_1_d_bits_sink;
  wire [31:0] TLBuffer_3_io_out_1_d_bits_data;
  wire  TLBuffer_3_io_out_1_d_bits_error;
  wire  TLBuffer_3_io_out_0_a_ready;
  wire  TLBuffer_3_io_out_0_a_valid;
  wire [2:0] TLBuffer_3_io_out_0_a_bits_opcode;
  wire [2:0] TLBuffer_3_io_out_0_a_bits_size;
  wire [4:0] TLBuffer_3_io_out_0_a_bits_source;
  wire [27:0] TLBuffer_3_io_out_0_a_bits_address;
  wire [3:0] TLBuffer_3_io_out_0_a_bits_mask;
  wire [31:0] TLBuffer_3_io_out_0_a_bits_data;
  wire  TLBuffer_3_io_out_0_d_ready;
  wire  TLBuffer_3_io_out_0_d_valid;
  wire [2:0] TLBuffer_3_io_out_0_d_bits_opcode;
  wire [1:0] TLBuffer_3_io_out_0_d_bits_param;
  wire [2:0] TLBuffer_3_io_out_0_d_bits_size;
  wire [4:0] TLBuffer_3_io_out_0_d_bits_source;
  wire  TLBuffer_3_io_out_0_d_bits_sink;
  wire [31:0] TLBuffer_3_io_out_0_d_bits_data;
  wire  TLBuffer_3_io_out_0_d_bits_error;
  wire  TLFragmenter_1_clock;
  wire  TLFragmenter_1_reset;
  wire  TLFragmenter_1_io_in_3_a_ready;
  wire  TLFragmenter_1_io_in_3_a_valid;
  wire [2:0] TLFragmenter_1_io_in_3_a_bits_opcode;
  wire [2:0] TLFragmenter_1_io_in_3_a_bits_size;
  wire [4:0] TLFragmenter_1_io_in_3_a_bits_source;
  wire [16:0] TLFragmenter_1_io_in_3_a_bits_address;
  wire [3:0] TLFragmenter_1_io_in_3_a_bits_mask;
  wire  TLFragmenter_1_io_in_3_d_ready;
  wire  TLFragmenter_1_io_in_3_d_valid;
  wire [2:0] TLFragmenter_1_io_in_3_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_in_3_d_bits_param;
  wire [2:0] TLFragmenter_1_io_in_3_d_bits_size;
  wire [4:0] TLFragmenter_1_io_in_3_d_bits_source;
  wire  TLFragmenter_1_io_in_3_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_in_3_d_bits_data;
  wire  TLFragmenter_1_io_in_3_d_bits_error;
  wire  TLFragmenter_1_io_in_2_a_ready;
  wire  TLFragmenter_1_io_in_2_a_valid;
  wire [2:0] TLFragmenter_1_io_in_2_a_bits_opcode;
  wire [2:0] TLFragmenter_1_io_in_2_a_bits_size;
  wire [4:0] TLFragmenter_1_io_in_2_a_bits_source;
  wire [11:0] TLFragmenter_1_io_in_2_a_bits_address;
  wire [3:0] TLFragmenter_1_io_in_2_a_bits_mask;
  wire [31:0] TLFragmenter_1_io_in_2_a_bits_data;
  wire  TLFragmenter_1_io_in_2_d_ready;
  wire  TLFragmenter_1_io_in_2_d_valid;
  wire [2:0] TLFragmenter_1_io_in_2_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_in_2_d_bits_param;
  wire [2:0] TLFragmenter_1_io_in_2_d_bits_size;
  wire [4:0] TLFragmenter_1_io_in_2_d_bits_source;
  wire  TLFragmenter_1_io_in_2_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_in_2_d_bits_data;
  wire  TLFragmenter_1_io_in_2_d_bits_error;
  wire  TLFragmenter_1_io_in_1_a_ready;
  wire  TLFragmenter_1_io_in_1_a_valid;
  wire [2:0] TLFragmenter_1_io_in_1_a_bits_opcode;
  wire [2:0] TLFragmenter_1_io_in_1_a_bits_size;
  wire [4:0] TLFragmenter_1_io_in_1_a_bits_source;
  wire [25:0] TLFragmenter_1_io_in_1_a_bits_address;
  wire [3:0] TLFragmenter_1_io_in_1_a_bits_mask;
  wire [31:0] TLFragmenter_1_io_in_1_a_bits_data;
  wire  TLFragmenter_1_io_in_1_d_ready;
  wire  TLFragmenter_1_io_in_1_d_valid;
  wire [2:0] TLFragmenter_1_io_in_1_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_in_1_d_bits_param;
  wire [2:0] TLFragmenter_1_io_in_1_d_bits_size;
  wire [4:0] TLFragmenter_1_io_in_1_d_bits_source;
  wire  TLFragmenter_1_io_in_1_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_in_1_d_bits_data;
  wire  TLFragmenter_1_io_in_1_d_bits_error;
  wire  TLFragmenter_1_io_in_0_a_ready;
  wire  TLFragmenter_1_io_in_0_a_valid;
  wire [2:0] TLFragmenter_1_io_in_0_a_bits_opcode;
  wire [2:0] TLFragmenter_1_io_in_0_a_bits_size;
  wire [4:0] TLFragmenter_1_io_in_0_a_bits_source;
  wire [27:0] TLFragmenter_1_io_in_0_a_bits_address;
  wire [3:0] TLFragmenter_1_io_in_0_a_bits_mask;
  wire [31:0] TLFragmenter_1_io_in_0_a_bits_data;
  wire  TLFragmenter_1_io_in_0_d_ready;
  wire  TLFragmenter_1_io_in_0_d_valid;
  wire [2:0] TLFragmenter_1_io_in_0_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_in_0_d_bits_param;
  wire [2:0] TLFragmenter_1_io_in_0_d_bits_size;
  wire [4:0] TLFragmenter_1_io_in_0_d_bits_source;
  wire  TLFragmenter_1_io_in_0_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_in_0_d_bits_data;
  wire  TLFragmenter_1_io_in_0_d_bits_error;
  wire  TLFragmenter_1_io_out_3_a_ready;
  wire  TLFragmenter_1_io_out_3_a_valid;
  wire [1:0] TLFragmenter_1_io_out_3_a_bits_size;
  wire [9:0] TLFragmenter_1_io_out_3_a_bits_source;
  wire [16:0] TLFragmenter_1_io_out_3_a_bits_address;
  wire  TLFragmenter_1_io_out_3_d_ready;
  wire  TLFragmenter_1_io_out_3_d_valid;
  wire [2:0] TLFragmenter_1_io_out_3_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_3_d_bits_param;
  wire [1:0] TLFragmenter_1_io_out_3_d_bits_size;
  wire [9:0] TLFragmenter_1_io_out_3_d_bits_source;
  wire  TLFragmenter_1_io_out_3_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_out_3_d_bits_data;
  wire  TLFragmenter_1_io_out_3_d_bits_error;
  wire  TLFragmenter_1_io_out_2_a_ready;
  wire  TLFragmenter_1_io_out_2_a_valid;
  wire [2:0] TLFragmenter_1_io_out_2_a_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_2_a_bits_size;
  wire [9:0] TLFragmenter_1_io_out_2_a_bits_source;
  wire [11:0] TLFragmenter_1_io_out_2_a_bits_address;
  wire [3:0] TLFragmenter_1_io_out_2_a_bits_mask;
  wire [31:0] TLFragmenter_1_io_out_2_a_bits_data;
  wire  TLFragmenter_1_io_out_2_d_ready;
  wire  TLFragmenter_1_io_out_2_d_valid;
  wire [2:0] TLFragmenter_1_io_out_2_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_2_d_bits_param;
  wire [1:0] TLFragmenter_1_io_out_2_d_bits_size;
  wire [9:0] TLFragmenter_1_io_out_2_d_bits_source;
  wire  TLFragmenter_1_io_out_2_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_out_2_d_bits_data;
  wire  TLFragmenter_1_io_out_2_d_bits_error;
  wire  TLFragmenter_1_io_out_1_a_ready;
  wire  TLFragmenter_1_io_out_1_a_valid;
  wire [2:0] TLFragmenter_1_io_out_1_a_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_1_a_bits_size;
  wire [9:0] TLFragmenter_1_io_out_1_a_bits_source;
  wire [25:0] TLFragmenter_1_io_out_1_a_bits_address;
  wire [3:0] TLFragmenter_1_io_out_1_a_bits_mask;
  wire [31:0] TLFragmenter_1_io_out_1_a_bits_data;
  wire  TLFragmenter_1_io_out_1_d_ready;
  wire  TLFragmenter_1_io_out_1_d_valid;
  wire [2:0] TLFragmenter_1_io_out_1_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_1_d_bits_param;
  wire [1:0] TLFragmenter_1_io_out_1_d_bits_size;
  wire [9:0] TLFragmenter_1_io_out_1_d_bits_source;
  wire  TLFragmenter_1_io_out_1_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_out_1_d_bits_data;
  wire  TLFragmenter_1_io_out_1_d_bits_error;
  wire  TLFragmenter_1_io_out_0_a_ready;
  wire  TLFragmenter_1_io_out_0_a_valid;
  wire [2:0] TLFragmenter_1_io_out_0_a_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_0_a_bits_size;
  wire [9:0] TLFragmenter_1_io_out_0_a_bits_source;
  wire [27:0] TLFragmenter_1_io_out_0_a_bits_address;
  wire [3:0] TLFragmenter_1_io_out_0_a_bits_mask;
  wire [31:0] TLFragmenter_1_io_out_0_a_bits_data;
  wire  TLFragmenter_1_io_out_0_d_ready;
  wire  TLFragmenter_1_io_out_0_d_valid;
  wire [2:0] TLFragmenter_1_io_out_0_d_bits_opcode;
  wire [1:0] TLFragmenter_1_io_out_0_d_bits_param;
  wire [1:0] TLFragmenter_1_io_out_0_d_bits_size;
  wire [9:0] TLFragmenter_1_io_out_0_d_bits_source;
  wire  TLFragmenter_1_io_out_0_d_bits_sink;
  wire [31:0] TLFragmenter_1_io_out_0_d_bits_data;
  wire  TLFragmenter_1_io_out_0_d_bits_error;
  wire  TLAtomicAutomata_clock;
  wire  TLAtomicAutomata_reset;
  wire  TLAtomicAutomata_io_in_0_a_ready;
  wire  TLAtomicAutomata_io_in_0_a_valid;
  wire [2:0] TLAtomicAutomata_io_in_0_a_bits_opcode;
  wire [2:0] TLAtomicAutomata_io_in_0_a_bits_param;
  wire [2:0] TLAtomicAutomata_io_in_0_a_bits_size;
  wire [4:0] TLAtomicAutomata_io_in_0_a_bits_source;
  wire [31:0] TLAtomicAutomata_io_in_0_a_bits_address;
  wire [3:0] TLAtomicAutomata_io_in_0_a_bits_mask;
  wire [31:0] TLAtomicAutomata_io_in_0_a_bits_data;
  wire  TLAtomicAutomata_io_in_0_d_ready;
  wire  TLAtomicAutomata_io_in_0_d_valid;
  wire [2:0] TLAtomicAutomata_io_in_0_d_bits_opcode;
  wire [1:0] TLAtomicAutomata_io_in_0_d_bits_param;
  wire [2:0] TLAtomicAutomata_io_in_0_d_bits_size;
  wire [4:0] TLAtomicAutomata_io_in_0_d_bits_source;
  wire  TLAtomicAutomata_io_in_0_d_bits_sink;
  wire [31:0] TLAtomicAutomata_io_in_0_d_bits_data;
  wire  TLAtomicAutomata_io_in_0_d_bits_error;
  wire  TLAtomicAutomata_io_out_0_a_ready;
  wire  TLAtomicAutomata_io_out_0_a_valid;
  wire [2:0] TLAtomicAutomata_io_out_0_a_bits_opcode;
  wire [2:0] TLAtomicAutomata_io_out_0_a_bits_param;
  wire [2:0] TLAtomicAutomata_io_out_0_a_bits_size;
  wire [4:0] TLAtomicAutomata_io_out_0_a_bits_source;
  wire [31:0] TLAtomicAutomata_io_out_0_a_bits_address;
  wire [3:0] TLAtomicAutomata_io_out_0_a_bits_mask;
  wire [31:0] TLAtomicAutomata_io_out_0_a_bits_data;
  wire  TLAtomicAutomata_io_out_0_d_ready;
  wire  TLAtomicAutomata_io_out_0_d_valid;
  wire [2:0] TLAtomicAutomata_io_out_0_d_bits_opcode;
  wire [1:0] TLAtomicAutomata_io_out_0_d_bits_param;
  wire [2:0] TLAtomicAutomata_io_out_0_d_bits_size;
  wire [4:0] TLAtomicAutomata_io_out_0_d_bits_source;
  wire  TLAtomicAutomata_io_out_0_d_bits_sink;
  wire [31:0] TLAtomicAutomata_io_out_0_d_bits_data;
  wire  TLAtomicAutomata_io_out_0_d_bits_error;
  wire  plic_clock;
  wire  plic_reset;
  wire  plic_io_tl_in_0_a_ready;
  wire  plic_io_tl_in_0_a_valid;
  wire [2:0] plic_io_tl_in_0_a_bits_opcode;
  wire [1:0] plic_io_tl_in_0_a_bits_size;
  wire [9:0] plic_io_tl_in_0_a_bits_source;
  wire [27:0] plic_io_tl_in_0_a_bits_address;
  wire [3:0] plic_io_tl_in_0_a_bits_mask;
  wire [31:0] plic_io_tl_in_0_a_bits_data;
  wire  plic_io_tl_in_0_d_ready;
  wire  plic_io_tl_in_0_d_valid;
  wire [2:0] plic_io_tl_in_0_d_bits_opcode;
  wire [1:0] plic_io_tl_in_0_d_bits_param;
  wire [1:0] plic_io_tl_in_0_d_bits_size;
  wire [9:0] plic_io_tl_in_0_d_bits_source;
  wire  plic_io_tl_in_0_d_bits_sink;
  wire [31:0] plic_io_tl_in_0_d_bits_data;
  wire  plic_io_tl_in_0_d_bits_error;
  wire  plic_io_devices_0_0;
  wire  plic_io_devices_0_1;
  wire  plic_io_harts_0_0;
  wire  clint_clock;
  wire  clint_reset;
  wire  clint_io_rtcTick;
  wire  clint_io_int_0_0;
  wire  clint_io_int_0_1;
  wire  clint_io_in_0_a_ready;
  wire  clint_io_in_0_a_valid;
  wire [2:0] clint_io_in_0_a_bits_opcode;
  wire [1:0] clint_io_in_0_a_bits_size;
  wire [9:0] clint_io_in_0_a_bits_source;
  wire [25:0] clint_io_in_0_a_bits_address;
  wire [3:0] clint_io_in_0_a_bits_mask;
  wire [31:0] clint_io_in_0_a_bits_data;
  wire  clint_io_in_0_d_ready;
  wire  clint_io_in_0_d_valid;
  wire [2:0] clint_io_in_0_d_bits_opcode;
  wire [1:0] clint_io_in_0_d_bits_param;
  wire [1:0] clint_io_in_0_d_bits_size;
  wire [9:0] clint_io_in_0_d_bits_source;
  wire  clint_io_in_0_d_bits_sink;
  wire [31:0] clint_io_in_0_d_bits_data;
  wire  clint_io_in_0_d_bits_error;
  wire  debug_1_clock;
  wire  debug_1_reset;
  wire  debug_1_io_debugInterrupts_0_0;
  wire  debug_1_io_in_0_a_ready;
  wire  debug_1_io_in_0_a_valid;
  wire [2:0] debug_1_io_in_0_a_bits_opcode;
  wire [1:0] debug_1_io_in_0_a_bits_size;
  wire [9:0] debug_1_io_in_0_a_bits_source;
  wire [11:0] debug_1_io_in_0_a_bits_address;
  wire [3:0] debug_1_io_in_0_a_bits_mask;
  wire [31:0] debug_1_io_in_0_a_bits_data;
  wire  debug_1_io_in_0_d_ready;
  wire  debug_1_io_in_0_d_valid;
  wire [2:0] debug_1_io_in_0_d_bits_opcode;
  wire [1:0] debug_1_io_in_0_d_bits_param;
  wire [1:0] debug_1_io_in_0_d_bits_size;
  wire [9:0] debug_1_io_in_0_d_bits_source;
  wire  debug_1_io_in_0_d_bits_sink;
  wire [31:0] debug_1_io_in_0_d_bits_data;
  wire  debug_1_io_in_0_d_bits_error;
  wire  debug_1_io_ctrl_debugUnavail_0;
  wire  debug_1_io_ctrl_ndreset;
  wire  debug_1_io_dmi_dmi_req_ready;
  wire  debug_1_io_dmi_dmi_req_valid;
  wire [6:0] debug_1_io_dmi_dmi_req_bits_addr;
  wire [31:0] debug_1_io_dmi_dmi_req_bits_data;
  wire [1:0] debug_1_io_dmi_dmi_req_bits_op;
  wire  debug_1_io_dmi_dmi_resp_ready;
  wire  debug_1_io_dmi_dmi_resp_valid;
  wire [31:0] debug_1_io_dmi_dmi_resp_bits_data;
  wire [1:0] debug_1_io_dmi_dmi_resp_bits_resp;
  wire  debug_1_io_dmi_dmiClock;
  wire  debug_1_io_dmi_dmiReset;
  wire  tile_clock;
  wire  tile_reset;
  wire  tile_io_master_0_a_ready;
  wire  tile_io_master_0_a_valid;
  wire [2:0] tile_io_master_0_a_bits_opcode;
  wire [2:0] tile_io_master_0_a_bits_param;
  wire [3:0] tile_io_master_0_a_bits_size;
  wire  tile_io_master_0_a_bits_source;
  wire [31:0] tile_io_master_0_a_bits_address;
  wire [3:0] tile_io_master_0_a_bits_mask;
  wire [31:0] tile_io_master_0_a_bits_data;
  wire  tile_io_master_0_d_ready;
  wire  tile_io_master_0_d_valid;
  wire [2:0] tile_io_master_0_d_bits_opcode;
  wire [3:0] tile_io_master_0_d_bits_size;
  wire  tile_io_master_0_d_bits_source;
  wire [31:0] tile_io_master_0_d_bits_data;
  wire  tile_io_master_0_d_bits_error;
  wire  tile_io_slave_0_a_ready;
  wire  tile_io_slave_0_a_valid;
  wire [2:0] tile_io_slave_0_a_bits_opcode;
  wire [2:0] tile_io_slave_0_a_bits_param;
  wire [2:0] tile_io_slave_0_a_bits_size;
  wire [4:0] tile_io_slave_0_a_bits_source;
  wire [31:0] tile_io_slave_0_a_bits_address;
  wire [3:0] tile_io_slave_0_a_bits_mask;
  wire [31:0] tile_io_slave_0_a_bits_data;
  wire  tile_io_slave_0_d_ready;
  wire  tile_io_slave_0_d_valid;
  wire [2:0] tile_io_slave_0_d_bits_opcode;
  wire [1:0] tile_io_slave_0_d_bits_param;
  wire [2:0] tile_io_slave_0_d_bits_size;
  wire [4:0] tile_io_slave_0_d_bits_source;
  wire  tile_io_slave_0_d_bits_sink;
  wire [31:0] tile_io_slave_0_d_bits_data;
  wire  tile_io_slave_0_d_bits_error;
  wire  tile_io_asyncInterrupts_0_0;
  wire  tile_io_periphInterrupts_0_0;
  wire  tile_io_periphInterrupts_0_1;
  wire  tile_io_periphInterrupts_0_2;
  wire  tile_io_hartid;
  wire [31:0] tile_io_resetVector;
  wire  TLBuffer_4_clock;
  wire  TLBuffer_4_reset;
  wire  TLBuffer_4_io_in_0_a_ready;
  wire  TLBuffer_4_io_in_0_a_valid;
  wire [2:0] TLBuffer_4_io_in_0_a_bits_opcode;
  wire [2:0] TLBuffer_4_io_in_0_a_bits_param;
  wire [3:0] TLBuffer_4_io_in_0_a_bits_size;
  wire  TLBuffer_4_io_in_0_a_bits_source;
  wire [31:0] TLBuffer_4_io_in_0_a_bits_address;
  wire [3:0] TLBuffer_4_io_in_0_a_bits_mask;
  wire [31:0] TLBuffer_4_io_in_0_a_bits_data;
  wire  TLBuffer_4_io_in_0_d_ready;
  wire  TLBuffer_4_io_in_0_d_valid;
  wire [2:0] TLBuffer_4_io_in_0_d_bits_opcode;
  wire [3:0] TLBuffer_4_io_in_0_d_bits_size;
  wire  TLBuffer_4_io_in_0_d_bits_source;
  wire [31:0] TLBuffer_4_io_in_0_d_bits_data;
  wire  TLBuffer_4_io_in_0_d_bits_error;
  wire  TLBuffer_4_io_out_0_a_ready;
  wire  TLBuffer_4_io_out_0_a_valid;
  wire [2:0] TLBuffer_4_io_out_0_a_bits_opcode;
  wire [2:0] TLBuffer_4_io_out_0_a_bits_param;
  wire [3:0] TLBuffer_4_io_out_0_a_bits_size;
  wire  TLBuffer_4_io_out_0_a_bits_source;
  wire [31:0] TLBuffer_4_io_out_0_a_bits_address;
  wire [3:0] TLBuffer_4_io_out_0_a_bits_mask;
  wire [31:0] TLBuffer_4_io_out_0_a_bits_data;
  wire  TLBuffer_4_io_out_0_d_ready;
  wire  TLBuffer_4_io_out_0_d_valid;
  wire [2:0] TLBuffer_4_io_out_0_d_bits_opcode;
  wire [3:0] TLBuffer_4_io_out_0_d_bits_size;
  wire  TLBuffer_4_io_out_0_d_bits_source;
  wire [31:0] TLBuffer_4_io_out_0_d_bits_data;
  wire  TLBuffer_4_io_out_0_d_bits_error;
  wire  IntXbar_1_io_in_0_0;
  wire  IntXbar_1_io_out_0_0;
  wire  IntXbar_2_io_in_1_0;
  wire  IntXbar_2_io_in_0_0;
  wire  IntXbar_2_io_in_0_1;
  wire  IntXbar_2_io_out_0_0;
  wire  IntXbar_2_io_out_0_1;
  wire  IntXbar_2_io_out_0_2;
  wire  IntXing_clock;
  wire  IntXing_io_in_0_0;
  wire  IntXing_io_in_0_1;
  wire  IntXing_io_out_0_0;
  wire  IntXing_io_out_0_1;
  wire  TLToAXI4_clock;
  wire  TLToAXI4_reset;
  wire  TLToAXI4_io_in_0_a_ready;
  wire  TLToAXI4_io_in_0_a_valid;
  wire [2:0] TLToAXI4_io_in_0_a_bits_opcode;
  wire [3:0] TLToAXI4_io_in_0_a_bits_size;
  wire [4:0] TLToAXI4_io_in_0_a_bits_source;
  wire [30:0] TLToAXI4_io_in_0_a_bits_address;
  wire [7:0] TLToAXI4_io_in_0_a_bits_mask;
  wire [63:0] TLToAXI4_io_in_0_a_bits_data;
  wire  TLToAXI4_io_in_0_d_ready;
  wire  TLToAXI4_io_in_0_d_valid;
  wire [2:0] TLToAXI4_io_in_0_d_bits_opcode;
  wire [1:0] TLToAXI4_io_in_0_d_bits_param;
  wire [3:0] TLToAXI4_io_in_0_d_bits_size;
  wire [4:0] TLToAXI4_io_in_0_d_bits_source;
  wire  TLToAXI4_io_in_0_d_bits_sink;
  wire [63:0] TLToAXI4_io_in_0_d_bits_data;
  wire  TLToAXI4_io_in_0_d_bits_error;
  wire  TLToAXI4_io_out_0_aw_ready;
  wire  TLToAXI4_io_out_0_aw_valid;
  wire [1:0] TLToAXI4_io_out_0_aw_bits_id;
  wire [30:0] TLToAXI4_io_out_0_aw_bits_addr;
  wire [7:0] TLToAXI4_io_out_0_aw_bits_len;
  wire [2:0] TLToAXI4_io_out_0_aw_bits_size;
  wire [1:0] TLToAXI4_io_out_0_aw_bits_burst;
  wire [11:0] TLToAXI4_io_out_0_aw_bits_user;
  wire  TLToAXI4_io_out_0_w_ready;
  wire  TLToAXI4_io_out_0_w_valid;
  wire [63:0] TLToAXI4_io_out_0_w_bits_data;
  wire [7:0] TLToAXI4_io_out_0_w_bits_strb;
  wire  TLToAXI4_io_out_0_w_bits_last;
  wire  TLToAXI4_io_out_0_b_ready;
  wire  TLToAXI4_io_out_0_b_valid;
  wire [1:0] TLToAXI4_io_out_0_b_bits_id;
  wire [1:0] TLToAXI4_io_out_0_b_bits_resp;
  wire [11:0] TLToAXI4_io_out_0_b_bits_user;
  wire  TLToAXI4_io_out_0_ar_ready;
  wire  TLToAXI4_io_out_0_ar_valid;
  wire [1:0] TLToAXI4_io_out_0_ar_bits_id;
  wire [30:0] TLToAXI4_io_out_0_ar_bits_addr;
  wire [7:0] TLToAXI4_io_out_0_ar_bits_len;
  wire [2:0] TLToAXI4_io_out_0_ar_bits_size;
  wire [1:0] TLToAXI4_io_out_0_ar_bits_burst;
  wire [11:0] TLToAXI4_io_out_0_ar_bits_user;
  wire  TLToAXI4_io_out_0_r_ready;
  wire  TLToAXI4_io_out_0_r_valid;
  wire [1:0] TLToAXI4_io_out_0_r_bits_id;
  wire [63:0] TLToAXI4_io_out_0_r_bits_data;
  wire [1:0] TLToAXI4_io_out_0_r_bits_resp;
  wire [11:0] TLToAXI4_io_out_0_r_bits_user;
  wire  TLToAXI4_io_out_0_r_bits_last;
  wire  AXI4IdIndexer_io_in_0_aw_ready;
  wire  AXI4IdIndexer_io_in_0_aw_valid;
  wire [1:0] AXI4IdIndexer_io_in_0_aw_bits_id;
  wire [30:0] AXI4IdIndexer_io_in_0_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_io_in_0_aw_bits_len;
  wire [2:0] AXI4IdIndexer_io_in_0_aw_bits_size;
  wire [1:0] AXI4IdIndexer_io_in_0_aw_bits_burst;
  wire [11:0] AXI4IdIndexer_io_in_0_aw_bits_user;
  wire  AXI4IdIndexer_io_in_0_w_ready;
  wire  AXI4IdIndexer_io_in_0_w_valid;
  wire [63:0] AXI4IdIndexer_io_in_0_w_bits_data;
  wire [7:0] AXI4IdIndexer_io_in_0_w_bits_strb;
  wire  AXI4IdIndexer_io_in_0_w_bits_last;
  wire  AXI4IdIndexer_io_in_0_b_ready;
  wire  AXI4IdIndexer_io_in_0_b_valid;
  wire [1:0] AXI4IdIndexer_io_in_0_b_bits_id;
  wire [1:0] AXI4IdIndexer_io_in_0_b_bits_resp;
  wire [11:0] AXI4IdIndexer_io_in_0_b_bits_user;
  wire  AXI4IdIndexer_io_in_0_ar_ready;
  wire  AXI4IdIndexer_io_in_0_ar_valid;
  wire [1:0] AXI4IdIndexer_io_in_0_ar_bits_id;
  wire [30:0] AXI4IdIndexer_io_in_0_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_io_in_0_ar_bits_len;
  wire [2:0] AXI4IdIndexer_io_in_0_ar_bits_size;
  wire [1:0] AXI4IdIndexer_io_in_0_ar_bits_burst;
  wire [11:0] AXI4IdIndexer_io_in_0_ar_bits_user;
  wire  AXI4IdIndexer_io_in_0_r_ready;
  wire  AXI4IdIndexer_io_in_0_r_valid;
  wire [1:0] AXI4IdIndexer_io_in_0_r_bits_id;
  wire [63:0] AXI4IdIndexer_io_in_0_r_bits_data;
  wire [1:0] AXI4IdIndexer_io_in_0_r_bits_resp;
  wire [11:0] AXI4IdIndexer_io_in_0_r_bits_user;
  wire  AXI4IdIndexer_io_in_0_r_bits_last;
  wire  AXI4IdIndexer_io_out_0_aw_ready;
  wire  AXI4IdIndexer_io_out_0_aw_valid;
  wire [3:0] AXI4IdIndexer_io_out_0_aw_bits_id;
  wire [30:0] AXI4IdIndexer_io_out_0_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_io_out_0_aw_bits_len;
  wire [2:0] AXI4IdIndexer_io_out_0_aw_bits_size;
  wire [1:0] AXI4IdIndexer_io_out_0_aw_bits_burst;
  wire [11:0] AXI4IdIndexer_io_out_0_aw_bits_user;
  wire  AXI4IdIndexer_io_out_0_w_ready;
  wire  AXI4IdIndexer_io_out_0_w_valid;
  wire [63:0] AXI4IdIndexer_io_out_0_w_bits_data;
  wire [7:0] AXI4IdIndexer_io_out_0_w_bits_strb;
  wire  AXI4IdIndexer_io_out_0_w_bits_last;
  wire  AXI4IdIndexer_io_out_0_b_ready;
  wire  AXI4IdIndexer_io_out_0_b_valid;
  wire [3:0] AXI4IdIndexer_io_out_0_b_bits_id;
  wire [1:0] AXI4IdIndexer_io_out_0_b_bits_resp;
  wire [11:0] AXI4IdIndexer_io_out_0_b_bits_user;
  wire  AXI4IdIndexer_io_out_0_ar_ready;
  wire  AXI4IdIndexer_io_out_0_ar_valid;
  wire [3:0] AXI4IdIndexer_io_out_0_ar_bits_id;
  wire [30:0] AXI4IdIndexer_io_out_0_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_io_out_0_ar_bits_len;
  wire [2:0] AXI4IdIndexer_io_out_0_ar_bits_size;
  wire [1:0] AXI4IdIndexer_io_out_0_ar_bits_burst;
  wire [11:0] AXI4IdIndexer_io_out_0_ar_bits_user;
  wire  AXI4IdIndexer_io_out_0_r_ready;
  wire  AXI4IdIndexer_io_out_0_r_valid;
  wire [3:0] AXI4IdIndexer_io_out_0_r_bits_id;
  wire [63:0] AXI4IdIndexer_io_out_0_r_bits_data;
  wire [1:0] AXI4IdIndexer_io_out_0_r_bits_resp;
  wire [11:0] AXI4IdIndexer_io_out_0_r_bits_user;
  wire  AXI4IdIndexer_io_out_0_r_bits_last;
  wire  AXI4Deinterleaver_clock;
  wire  AXI4Deinterleaver_reset;
  wire  AXI4Deinterleaver_io_in_0_aw_ready;
  wire  AXI4Deinterleaver_io_in_0_aw_valid;
  wire [3:0] AXI4Deinterleaver_io_in_0_aw_bits_id;
  wire [30:0] AXI4Deinterleaver_io_in_0_aw_bits_addr;
  wire [7:0] AXI4Deinterleaver_io_in_0_aw_bits_len;
  wire [2:0] AXI4Deinterleaver_io_in_0_aw_bits_size;
  wire [1:0] AXI4Deinterleaver_io_in_0_aw_bits_burst;
  wire [11:0] AXI4Deinterleaver_io_in_0_aw_bits_user;
  wire  AXI4Deinterleaver_io_in_0_w_ready;
  wire  AXI4Deinterleaver_io_in_0_w_valid;
  wire [63:0] AXI4Deinterleaver_io_in_0_w_bits_data;
  wire [7:0] AXI4Deinterleaver_io_in_0_w_bits_strb;
  wire  AXI4Deinterleaver_io_in_0_w_bits_last;
  wire  AXI4Deinterleaver_io_in_0_b_ready;
  wire  AXI4Deinterleaver_io_in_0_b_valid;
  wire [3:0] AXI4Deinterleaver_io_in_0_b_bits_id;
  wire [1:0] AXI4Deinterleaver_io_in_0_b_bits_resp;
  wire [11:0] AXI4Deinterleaver_io_in_0_b_bits_user;
  wire  AXI4Deinterleaver_io_in_0_ar_ready;
  wire  AXI4Deinterleaver_io_in_0_ar_valid;
  wire [3:0] AXI4Deinterleaver_io_in_0_ar_bits_id;
  wire [30:0] AXI4Deinterleaver_io_in_0_ar_bits_addr;
  wire [7:0] AXI4Deinterleaver_io_in_0_ar_bits_len;
  wire [2:0] AXI4Deinterleaver_io_in_0_ar_bits_size;
  wire [1:0] AXI4Deinterleaver_io_in_0_ar_bits_burst;
  wire [11:0] AXI4Deinterleaver_io_in_0_ar_bits_user;
  wire  AXI4Deinterleaver_io_in_0_r_ready;
  wire  AXI4Deinterleaver_io_in_0_r_valid;
  wire [3:0] AXI4Deinterleaver_io_in_0_r_bits_id;
  wire [63:0] AXI4Deinterleaver_io_in_0_r_bits_data;
  wire [1:0] AXI4Deinterleaver_io_in_0_r_bits_resp;
  wire [11:0] AXI4Deinterleaver_io_in_0_r_bits_user;
  wire  AXI4Deinterleaver_io_in_0_r_bits_last;
  wire  AXI4Deinterleaver_io_out_0_aw_ready;
  wire  AXI4Deinterleaver_io_out_0_aw_valid;
  wire [3:0] AXI4Deinterleaver_io_out_0_aw_bits_id;
  wire [30:0] AXI4Deinterleaver_io_out_0_aw_bits_addr;
  wire [7:0] AXI4Deinterleaver_io_out_0_aw_bits_len;
  wire [2:0] AXI4Deinterleaver_io_out_0_aw_bits_size;
  wire [1:0] AXI4Deinterleaver_io_out_0_aw_bits_burst;
  wire [11:0] AXI4Deinterleaver_io_out_0_aw_bits_user;
  wire  AXI4Deinterleaver_io_out_0_w_ready;
  wire  AXI4Deinterleaver_io_out_0_w_valid;
  wire [63:0] AXI4Deinterleaver_io_out_0_w_bits_data;
  wire [7:0] AXI4Deinterleaver_io_out_0_w_bits_strb;
  wire  AXI4Deinterleaver_io_out_0_w_bits_last;
  wire  AXI4Deinterleaver_io_out_0_b_ready;
  wire  AXI4Deinterleaver_io_out_0_b_valid;
  wire [3:0] AXI4Deinterleaver_io_out_0_b_bits_id;
  wire [1:0] AXI4Deinterleaver_io_out_0_b_bits_resp;
  wire [11:0] AXI4Deinterleaver_io_out_0_b_bits_user;
  wire  AXI4Deinterleaver_io_out_0_ar_ready;
  wire  AXI4Deinterleaver_io_out_0_ar_valid;
  wire [3:0] AXI4Deinterleaver_io_out_0_ar_bits_id;
  wire [30:0] AXI4Deinterleaver_io_out_0_ar_bits_addr;
  wire [7:0] AXI4Deinterleaver_io_out_0_ar_bits_len;
  wire [2:0] AXI4Deinterleaver_io_out_0_ar_bits_size;
  wire [1:0] AXI4Deinterleaver_io_out_0_ar_bits_burst;
  wire [11:0] AXI4Deinterleaver_io_out_0_ar_bits_user;
  wire  AXI4Deinterleaver_io_out_0_r_ready;
  wire  AXI4Deinterleaver_io_out_0_r_valid;
  wire [3:0] AXI4Deinterleaver_io_out_0_r_bits_id;
  wire [63:0] AXI4Deinterleaver_io_out_0_r_bits_data;
  wire [1:0] AXI4Deinterleaver_io_out_0_r_bits_resp;
  wire [11:0] AXI4Deinterleaver_io_out_0_r_bits_user;
  wire  AXI4Deinterleaver_io_out_0_r_bits_last;
  wire  AXI4UserYanker_clock;
  wire  AXI4UserYanker_reset;
  wire  AXI4UserYanker_io_in_0_aw_ready;
  wire  AXI4UserYanker_io_in_0_aw_valid;
  wire [3:0] AXI4UserYanker_io_in_0_aw_bits_id;
  wire [30:0] AXI4UserYanker_io_in_0_aw_bits_addr;
  wire [7:0] AXI4UserYanker_io_in_0_aw_bits_len;
  wire [2:0] AXI4UserYanker_io_in_0_aw_bits_size;
  wire [1:0] AXI4UserYanker_io_in_0_aw_bits_burst;
  wire [11:0] AXI4UserYanker_io_in_0_aw_bits_user;
  wire  AXI4UserYanker_io_in_0_w_ready;
  wire  AXI4UserYanker_io_in_0_w_valid;
  wire [63:0] AXI4UserYanker_io_in_0_w_bits_data;
  wire [7:0] AXI4UserYanker_io_in_0_w_bits_strb;
  wire  AXI4UserYanker_io_in_0_w_bits_last;
  wire  AXI4UserYanker_io_in_0_b_ready;
  wire  AXI4UserYanker_io_in_0_b_valid;
  wire [3:0] AXI4UserYanker_io_in_0_b_bits_id;
  wire [1:0] AXI4UserYanker_io_in_0_b_bits_resp;
  wire [11:0] AXI4UserYanker_io_in_0_b_bits_user;
  wire  AXI4UserYanker_io_in_0_ar_ready;
  wire  AXI4UserYanker_io_in_0_ar_valid;
  wire [3:0] AXI4UserYanker_io_in_0_ar_bits_id;
  wire [30:0] AXI4UserYanker_io_in_0_ar_bits_addr;
  wire [7:0] AXI4UserYanker_io_in_0_ar_bits_len;
  wire [2:0] AXI4UserYanker_io_in_0_ar_bits_size;
  wire [1:0] AXI4UserYanker_io_in_0_ar_bits_burst;
  wire [11:0] AXI4UserYanker_io_in_0_ar_bits_user;
  wire  AXI4UserYanker_io_in_0_r_ready;
  wire  AXI4UserYanker_io_in_0_r_valid;
  wire [3:0] AXI4UserYanker_io_in_0_r_bits_id;
  wire [63:0] AXI4UserYanker_io_in_0_r_bits_data;
  wire [1:0] AXI4UserYanker_io_in_0_r_bits_resp;
  wire [11:0] AXI4UserYanker_io_in_0_r_bits_user;
  wire  AXI4UserYanker_io_in_0_r_bits_last;
  wire  AXI4UserYanker_io_out_0_aw_ready;
  wire  AXI4UserYanker_io_out_0_aw_valid;
  wire [3:0] AXI4UserYanker_io_out_0_aw_bits_id;
  wire [30:0] AXI4UserYanker_io_out_0_aw_bits_addr;
  wire [7:0] AXI4UserYanker_io_out_0_aw_bits_len;
  wire [2:0] AXI4UserYanker_io_out_0_aw_bits_size;
  wire [1:0] AXI4UserYanker_io_out_0_aw_bits_burst;
  wire  AXI4UserYanker_io_out_0_w_ready;
  wire  AXI4UserYanker_io_out_0_w_valid;
  wire [63:0] AXI4UserYanker_io_out_0_w_bits_data;
  wire [7:0] AXI4UserYanker_io_out_0_w_bits_strb;
  wire  AXI4UserYanker_io_out_0_w_bits_last;
  wire  AXI4UserYanker_io_out_0_b_ready;
  wire  AXI4UserYanker_io_out_0_b_valid;
  wire [3:0] AXI4UserYanker_io_out_0_b_bits_id;
  wire [1:0] AXI4UserYanker_io_out_0_b_bits_resp;
  wire  AXI4UserYanker_io_out_0_ar_ready;
  wire  AXI4UserYanker_io_out_0_ar_valid;
  wire [3:0] AXI4UserYanker_io_out_0_ar_bits_id;
  wire [30:0] AXI4UserYanker_io_out_0_ar_bits_addr;
  wire [7:0] AXI4UserYanker_io_out_0_ar_bits_len;
  wire [2:0] AXI4UserYanker_io_out_0_ar_bits_size;
  wire [1:0] AXI4UserYanker_io_out_0_ar_bits_burst;
  wire  AXI4UserYanker_io_out_0_r_ready;
  wire  AXI4UserYanker_io_out_0_r_valid;
  wire [3:0] AXI4UserYanker_io_out_0_r_bits_id;
  wire [63:0] AXI4UserYanker_io_out_0_r_bits_data;
  wire [1:0] AXI4UserYanker_io_out_0_r_bits_resp;
  wire  AXI4UserYanker_io_out_0_r_bits_last;
  wire  AXI4Buffer_clock;
  wire  AXI4Buffer_reset;
  wire  AXI4Buffer_io_in_0_aw_ready;
  wire  AXI4Buffer_io_in_0_aw_valid;
  wire [3:0] AXI4Buffer_io_in_0_aw_bits_id;
  wire [30:0] AXI4Buffer_io_in_0_aw_bits_addr;
  wire [7:0] AXI4Buffer_io_in_0_aw_bits_len;
  wire [2:0] AXI4Buffer_io_in_0_aw_bits_size;
  wire [1:0] AXI4Buffer_io_in_0_aw_bits_burst;
  wire  AXI4Buffer_io_in_0_w_ready;
  wire  AXI4Buffer_io_in_0_w_valid;
  wire [63:0] AXI4Buffer_io_in_0_w_bits_data;
  wire [7:0] AXI4Buffer_io_in_0_w_bits_strb;
  wire  AXI4Buffer_io_in_0_w_bits_last;
  wire  AXI4Buffer_io_in_0_b_ready;
  wire  AXI4Buffer_io_in_0_b_valid;
  wire [3:0] AXI4Buffer_io_in_0_b_bits_id;
  wire [1:0] AXI4Buffer_io_in_0_b_bits_resp;
  wire  AXI4Buffer_io_in_0_ar_ready;
  wire  AXI4Buffer_io_in_0_ar_valid;
  wire [3:0] AXI4Buffer_io_in_0_ar_bits_id;
  wire [30:0] AXI4Buffer_io_in_0_ar_bits_addr;
  wire [7:0] AXI4Buffer_io_in_0_ar_bits_len;
  wire [2:0] AXI4Buffer_io_in_0_ar_bits_size;
  wire [1:0] AXI4Buffer_io_in_0_ar_bits_burst;
  wire  AXI4Buffer_io_in_0_r_ready;
  wire  AXI4Buffer_io_in_0_r_valid;
  wire [3:0] AXI4Buffer_io_in_0_r_bits_id;
  wire [63:0] AXI4Buffer_io_in_0_r_bits_data;
  wire [1:0] AXI4Buffer_io_in_0_r_bits_resp;
  wire  AXI4Buffer_io_in_0_r_bits_last;
  wire  AXI4Buffer_io_out_0_aw_ready;
  wire  AXI4Buffer_io_out_0_aw_valid;
  wire [3:0] AXI4Buffer_io_out_0_aw_bits_id;
  wire [30:0] AXI4Buffer_io_out_0_aw_bits_addr;
  wire [7:0] AXI4Buffer_io_out_0_aw_bits_len;
  wire [2:0] AXI4Buffer_io_out_0_aw_bits_size;
  wire [1:0] AXI4Buffer_io_out_0_aw_bits_burst;
  wire  AXI4Buffer_io_out_0_w_ready;
  wire  AXI4Buffer_io_out_0_w_valid;
  wire [63:0] AXI4Buffer_io_out_0_w_bits_data;
  wire [7:0] AXI4Buffer_io_out_0_w_bits_strb;
  wire  AXI4Buffer_io_out_0_w_bits_last;
  wire  AXI4Buffer_io_out_0_b_ready;
  wire  AXI4Buffer_io_out_0_b_valid;
  wire [3:0] AXI4Buffer_io_out_0_b_bits_id;
  wire [1:0] AXI4Buffer_io_out_0_b_bits_resp;
  wire  AXI4Buffer_io_out_0_ar_ready;
  wire  AXI4Buffer_io_out_0_ar_valid;
  wire [3:0] AXI4Buffer_io_out_0_ar_bits_id;
  wire [30:0] AXI4Buffer_io_out_0_ar_bits_addr;
  wire [7:0] AXI4Buffer_io_out_0_ar_bits_len;
  wire [2:0] AXI4Buffer_io_out_0_ar_bits_size;
  wire [1:0] AXI4Buffer_io_out_0_ar_bits_burst;
  wire  AXI4Buffer_io_out_0_r_ready;
  wire  AXI4Buffer_io_out_0_r_valid;
  wire [3:0] AXI4Buffer_io_out_0_r_bits_id;
  wire [63:0] AXI4Buffer_io_out_0_r_bits_data;
  wire [1:0] AXI4Buffer_io_out_0_r_bits_resp;
  wire  AXI4Buffer_io_out_0_r_bits_last;
  wire  TLBuffer_5_clock;
  wire  TLBuffer_5_reset;
  wire  TLBuffer_5_io_in_0_a_ready;
  wire  TLBuffer_5_io_in_0_a_valid;
  wire [2:0] TLBuffer_5_io_in_0_a_bits_opcode;
  wire [2:0] TLBuffer_5_io_in_0_a_bits_param;
  wire [3:0] TLBuffer_5_io_in_0_a_bits_size;
  wire [3:0] TLBuffer_5_io_in_0_a_bits_source;
  wire [31:0] TLBuffer_5_io_in_0_a_bits_address;
  wire [3:0] TLBuffer_5_io_in_0_a_bits_mask;
  wire [31:0] TLBuffer_5_io_in_0_a_bits_data;
  wire  TLBuffer_5_io_in_0_d_ready;
  wire  TLBuffer_5_io_in_0_d_valid;
  wire [2:0] TLBuffer_5_io_in_0_d_bits_opcode;
  wire [3:0] TLBuffer_5_io_in_0_d_bits_size;
  wire [3:0] TLBuffer_5_io_in_0_d_bits_source;
  wire  TLBuffer_5_io_out_0_a_ready;
  wire  TLBuffer_5_io_out_0_a_valid;
  wire [2:0] TLBuffer_5_io_out_0_a_bits_opcode;
  wire [2:0] TLBuffer_5_io_out_0_a_bits_param;
  wire [3:0] TLBuffer_5_io_out_0_a_bits_size;
  wire [3:0] TLBuffer_5_io_out_0_a_bits_source;
  wire [31:0] TLBuffer_5_io_out_0_a_bits_address;
  wire [3:0] TLBuffer_5_io_out_0_a_bits_mask;
  wire [31:0] TLBuffer_5_io_out_0_a_bits_data;
  wire  TLBuffer_5_io_out_0_d_ready;
  wire  TLBuffer_5_io_out_0_d_valid;
  wire [2:0] TLBuffer_5_io_out_0_d_bits_opcode;
  wire [3:0] TLBuffer_5_io_out_0_d_bits_size;
  wire [3:0] TLBuffer_5_io_out_0_d_bits_source;
  wire  AXI4IdIndexer_1_io_in_0_aw_valid;
  wire [7:0] AXI4IdIndexer_1_io_in_0_aw_bits_id;
  wire [31:0] AXI4IdIndexer_1_io_in_0_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_1_io_in_0_aw_bits_len;
  wire [2:0] AXI4IdIndexer_1_io_in_0_aw_bits_size;
  wire [1:0] AXI4IdIndexer_1_io_in_0_aw_bits_burst;
  wire  AXI4IdIndexer_1_io_in_0_w_valid;
  wire [63:0] AXI4IdIndexer_1_io_in_0_w_bits_data;
  wire [7:0] AXI4IdIndexer_1_io_in_0_w_bits_strb;
  wire  AXI4IdIndexer_1_io_in_0_w_bits_last;
  wire  AXI4IdIndexer_1_io_in_0_b_ready;
  wire  AXI4IdIndexer_1_io_in_0_ar_valid;
  wire [7:0] AXI4IdIndexer_1_io_in_0_ar_bits_id;
  wire [31:0] AXI4IdIndexer_1_io_in_0_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_1_io_in_0_ar_bits_len;
  wire [2:0] AXI4IdIndexer_1_io_in_0_ar_bits_size;
  wire [1:0] AXI4IdIndexer_1_io_in_0_ar_bits_burst;
  wire  AXI4IdIndexer_1_io_in_0_r_ready;
  wire  AXI4IdIndexer_1_io_out_0_aw_valid;
  wire  AXI4IdIndexer_1_io_out_0_aw_bits_id;
  wire [31:0] AXI4IdIndexer_1_io_out_0_aw_bits_addr;
  wire [7:0] AXI4IdIndexer_1_io_out_0_aw_bits_len;
  wire [2:0] AXI4IdIndexer_1_io_out_0_aw_bits_size;
  wire [1:0] AXI4IdIndexer_1_io_out_0_aw_bits_burst;
  wire [6:0] AXI4IdIndexer_1_io_out_0_aw_bits_user;
  wire  AXI4IdIndexer_1_io_out_0_w_valid;
  wire [63:0] AXI4IdIndexer_1_io_out_0_w_bits_data;
  wire [7:0] AXI4IdIndexer_1_io_out_0_w_bits_strb;
  wire  AXI4IdIndexer_1_io_out_0_w_bits_last;
  wire  AXI4IdIndexer_1_io_out_0_b_ready;
  wire  AXI4IdIndexer_1_io_out_0_ar_valid;
  wire  AXI4IdIndexer_1_io_out_0_ar_bits_id;
  wire [31:0] AXI4IdIndexer_1_io_out_0_ar_bits_addr;
  wire [7:0] AXI4IdIndexer_1_io_out_0_ar_bits_len;
  wire [2:0] AXI4IdIndexer_1_io_out_0_ar_bits_size;
  wire [1:0] AXI4IdIndexer_1_io_out_0_ar_bits_burst;
  wire [6:0] AXI4IdIndexer_1_io_out_0_ar_bits_user;
  wire  AXI4IdIndexer_1_io_out_0_r_ready;
  wire  AXI4Fragmenter_clock;
  wire  AXI4Fragmenter_reset;
  wire  AXI4Fragmenter_io_in_0_aw_valid;
  wire  AXI4Fragmenter_io_in_0_aw_bits_id;
  wire [31:0] AXI4Fragmenter_io_in_0_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_io_in_0_aw_bits_len;
  wire [2:0] AXI4Fragmenter_io_in_0_aw_bits_size;
  wire [1:0] AXI4Fragmenter_io_in_0_aw_bits_burst;
  wire [6:0] AXI4Fragmenter_io_in_0_aw_bits_user;
  wire  AXI4Fragmenter_io_in_0_w_valid;
  wire [63:0] AXI4Fragmenter_io_in_0_w_bits_data;
  wire [7:0] AXI4Fragmenter_io_in_0_w_bits_strb;
  wire  AXI4Fragmenter_io_in_0_w_bits_last;
  wire  AXI4Fragmenter_io_in_0_b_ready;
  wire  AXI4Fragmenter_io_in_0_ar_valid;
  wire  AXI4Fragmenter_io_in_0_ar_bits_id;
  wire [31:0] AXI4Fragmenter_io_in_0_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_io_in_0_ar_bits_len;
  wire [2:0] AXI4Fragmenter_io_in_0_ar_bits_size;
  wire [1:0] AXI4Fragmenter_io_in_0_ar_bits_burst;
  wire [6:0] AXI4Fragmenter_io_in_0_ar_bits_user;
  wire  AXI4Fragmenter_io_in_0_r_ready;
  wire  AXI4Fragmenter_io_out_0_aw_ready;
  wire  AXI4Fragmenter_io_out_0_aw_valid;
  wire  AXI4Fragmenter_io_out_0_aw_bits_id;
  wire [31:0] AXI4Fragmenter_io_out_0_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_io_out_0_aw_bits_len;
  wire [2:0] AXI4Fragmenter_io_out_0_aw_bits_size;
  wire [7:0] AXI4Fragmenter_io_out_0_aw_bits_user;
  wire  AXI4Fragmenter_io_out_0_w_ready;
  wire  AXI4Fragmenter_io_out_0_w_valid;
  wire [63:0] AXI4Fragmenter_io_out_0_w_bits_data;
  wire [7:0] AXI4Fragmenter_io_out_0_w_bits_strb;
  wire  AXI4Fragmenter_io_out_0_w_bits_last;
  wire  AXI4Fragmenter_io_out_0_b_ready;
  wire [7:0] AXI4Fragmenter_io_out_0_b_bits_user;
  wire  AXI4Fragmenter_io_out_0_ar_ready;
  wire  AXI4Fragmenter_io_out_0_ar_valid;
  wire  AXI4Fragmenter_io_out_0_ar_bits_id;
  wire [31:0] AXI4Fragmenter_io_out_0_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_io_out_0_ar_bits_len;
  wire [2:0] AXI4Fragmenter_io_out_0_ar_bits_size;
  wire [7:0] AXI4Fragmenter_io_out_0_ar_bits_user;
  wire  AXI4Fragmenter_io_out_0_r_ready;
  wire  AXI4UserYanker_1_clock;
  wire  AXI4UserYanker_1_reset;
  wire  AXI4UserYanker_1_io_in_0_aw_ready;
  wire  AXI4UserYanker_1_io_in_0_aw_valid;
  wire  AXI4UserYanker_1_io_in_0_aw_bits_id;
  wire [31:0] AXI4UserYanker_1_io_in_0_aw_bits_addr;
  wire [7:0] AXI4UserYanker_1_io_in_0_aw_bits_len;
  wire [2:0] AXI4UserYanker_1_io_in_0_aw_bits_size;
  wire [7:0] AXI4UserYanker_1_io_in_0_aw_bits_user;
  wire  AXI4UserYanker_1_io_in_0_w_ready;
  wire  AXI4UserYanker_1_io_in_0_w_valid;
  wire [63:0] AXI4UserYanker_1_io_in_0_w_bits_data;
  wire [7:0] AXI4UserYanker_1_io_in_0_w_bits_strb;
  wire  AXI4UserYanker_1_io_in_0_w_bits_last;
  wire  AXI4UserYanker_1_io_in_0_b_ready;
  wire [7:0] AXI4UserYanker_1_io_in_0_b_bits_user;
  wire  AXI4UserYanker_1_io_in_0_ar_ready;
  wire  AXI4UserYanker_1_io_in_0_ar_valid;
  wire  AXI4UserYanker_1_io_in_0_ar_bits_id;
  wire [31:0] AXI4UserYanker_1_io_in_0_ar_bits_addr;
  wire [7:0] AXI4UserYanker_1_io_in_0_ar_bits_len;
  wire [2:0] AXI4UserYanker_1_io_in_0_ar_bits_size;
  wire [7:0] AXI4UserYanker_1_io_in_0_ar_bits_user;
  wire  AXI4UserYanker_1_io_in_0_r_ready;
  wire  AXI4UserYanker_1_io_out_0_aw_ready;
  wire  AXI4UserYanker_1_io_out_0_aw_valid;
  wire  AXI4UserYanker_1_io_out_0_aw_bits_id;
  wire [31:0] AXI4UserYanker_1_io_out_0_aw_bits_addr;
  wire [7:0] AXI4UserYanker_1_io_out_0_aw_bits_len;
  wire [2:0] AXI4UserYanker_1_io_out_0_aw_bits_size;
  wire  AXI4UserYanker_1_io_out_0_w_ready;
  wire  AXI4UserYanker_1_io_out_0_w_valid;
  wire [63:0] AXI4UserYanker_1_io_out_0_w_bits_data;
  wire [7:0] AXI4UserYanker_1_io_out_0_w_bits_strb;
  wire  AXI4UserYanker_1_io_out_0_w_bits_last;
  wire  AXI4UserYanker_1_io_out_0_b_ready;
  wire  AXI4UserYanker_1_io_out_0_b_valid;
  wire  AXI4UserYanker_1_io_out_0_b_bits_id;
  wire  AXI4UserYanker_1_io_out_0_ar_ready;
  wire  AXI4UserYanker_1_io_out_0_ar_valid;
  wire  AXI4UserYanker_1_io_out_0_ar_bits_id;
  wire [31:0] AXI4UserYanker_1_io_out_0_ar_bits_addr;
  wire [7:0] AXI4UserYanker_1_io_out_0_ar_bits_len;
  wire [2:0] AXI4UserYanker_1_io_out_0_ar_bits_size;
  wire  AXI4UserYanker_1_io_out_0_r_ready;
  wire  AXI4UserYanker_1_io_out_0_r_valid;
  wire  AXI4UserYanker_1_io_out_0_r_bits_id;
  wire  AXI4UserYanker_1_io_out_0_r_bits_last;
  wire  AXI4ToTL_clock;
  wire  AXI4ToTL_reset;
  wire  AXI4ToTL_io_in_0_aw_ready;
  wire  AXI4ToTL_io_in_0_aw_valid;
  wire  AXI4ToTL_io_in_0_aw_bits_id;
  wire [31:0] AXI4ToTL_io_in_0_aw_bits_addr;
  wire [7:0] AXI4ToTL_io_in_0_aw_bits_len;
  wire [2:0] AXI4ToTL_io_in_0_aw_bits_size;
  wire  AXI4ToTL_io_in_0_w_ready;
  wire  AXI4ToTL_io_in_0_w_valid;
  wire [63:0] AXI4ToTL_io_in_0_w_bits_data;
  wire [7:0] AXI4ToTL_io_in_0_w_bits_strb;
  wire  AXI4ToTL_io_in_0_w_bits_last;
  wire  AXI4ToTL_io_in_0_b_ready;
  wire  AXI4ToTL_io_in_0_b_valid;
  wire  AXI4ToTL_io_in_0_b_bits_id;
  wire  AXI4ToTL_io_in_0_ar_ready;
  wire  AXI4ToTL_io_in_0_ar_valid;
  wire  AXI4ToTL_io_in_0_ar_bits_id;
  wire [31:0] AXI4ToTL_io_in_0_ar_bits_addr;
  wire [7:0] AXI4ToTL_io_in_0_ar_bits_len;
  wire [2:0] AXI4ToTL_io_in_0_ar_bits_size;
  wire  AXI4ToTL_io_in_0_r_ready;
  wire  AXI4ToTL_io_in_0_r_valid;
  wire  AXI4ToTL_io_in_0_r_bits_id;
  wire  AXI4ToTL_io_in_0_r_bits_last;
  wire  AXI4ToTL_io_out_0_a_ready;
  wire  AXI4ToTL_io_out_0_a_valid;
  wire [2:0] AXI4ToTL_io_out_0_a_bits_opcode;
  wire [2:0] AXI4ToTL_io_out_0_a_bits_param;
  wire [3:0] AXI4ToTL_io_out_0_a_bits_size;
  wire [3:0] AXI4ToTL_io_out_0_a_bits_source;
  wire [31:0] AXI4ToTL_io_out_0_a_bits_address;
  wire [7:0] AXI4ToTL_io_out_0_a_bits_mask;
  wire [63:0] AXI4ToTL_io_out_0_a_bits_data;
  wire  AXI4ToTL_io_out_0_d_ready;
  wire  AXI4ToTL_io_out_0_d_valid;
  wire [2:0] AXI4ToTL_io_out_0_d_bits_opcode;
  wire [3:0] AXI4ToTL_io_out_0_d_bits_size;
  wire [3:0] AXI4ToTL_io_out_0_d_bits_source;
  wire  TLWidthWidget_2_clock;
  wire  TLWidthWidget_2_reset;
  wire  TLWidthWidget_2_io_in_0_a_ready;
  wire  TLWidthWidget_2_io_in_0_a_valid;
  wire [2:0] TLWidthWidget_2_io_in_0_a_bits_opcode;
  wire [2:0] TLWidthWidget_2_io_in_0_a_bits_param;
  wire [3:0] TLWidthWidget_2_io_in_0_a_bits_size;
  wire [3:0] TLWidthWidget_2_io_in_0_a_bits_source;
  wire [31:0] TLWidthWidget_2_io_in_0_a_bits_address;
  wire [7:0] TLWidthWidget_2_io_in_0_a_bits_mask;
  wire [63:0] TLWidthWidget_2_io_in_0_a_bits_data;
  wire  TLWidthWidget_2_io_in_0_d_ready;
  wire  TLWidthWidget_2_io_in_0_d_valid;
  wire [2:0] TLWidthWidget_2_io_in_0_d_bits_opcode;
  wire [3:0] TLWidthWidget_2_io_in_0_d_bits_size;
  wire [3:0] TLWidthWidget_2_io_in_0_d_bits_source;
  wire  TLWidthWidget_2_io_out_0_a_ready;
  wire  TLWidthWidget_2_io_out_0_a_valid;
  wire [2:0] TLWidthWidget_2_io_out_0_a_bits_opcode;
  wire [2:0] TLWidthWidget_2_io_out_0_a_bits_param;
  wire [3:0] TLWidthWidget_2_io_out_0_a_bits_size;
  wire [3:0] TLWidthWidget_2_io_out_0_a_bits_source;
  wire [31:0] TLWidthWidget_2_io_out_0_a_bits_address;
  wire [3:0] TLWidthWidget_2_io_out_0_a_bits_mask;
  wire [31:0] TLWidthWidget_2_io_out_0_a_bits_data;
  wire  TLWidthWidget_2_io_out_0_d_ready;
  wire  TLWidthWidget_2_io_out_0_d_valid;
  wire [2:0] TLWidthWidget_2_io_out_0_d_bits_opcode;
  wire [3:0] TLWidthWidget_2_io_out_0_d_bits_size;
  wire [3:0] TLWidthWidget_2_io_out_0_d_bits_source;
  wire  bootrom_io_in_0_a_ready;
  wire  bootrom_io_in_0_a_valid;
  wire [1:0] bootrom_io_in_0_a_bits_size;
  wire [9:0] bootrom_io_in_0_a_bits_source;
  wire [16:0] bootrom_io_in_0_a_bits_address;
  wire  bootrom_io_in_0_d_ready;
  wire  bootrom_io_in_0_d_valid;
  wire [2:0] bootrom_io_in_0_d_bits_opcode;
  wire [1:0] bootrom_io_in_0_d_bits_param;
  wire [1:0] bootrom_io_in_0_d_bits_size;
  wire [9:0] bootrom_io_in_0_d_bits_source;
  wire  bootrom_io_in_0_d_bits_sink;
  wire [31:0] bootrom_io_in_0_d_bits_data;
  wire  bootrom_io_in_0_d_bits_error;
  wire  error_clock;
  wire  error_reset;
  wire  error_io_in_0_a_ready;
  wire  error_io_in_0_a_valid;
  wire [2:0] error_io_in_0_a_bits_opcode;
  wire [3:0] error_io_in_0_a_bits_size;
  wire [4:0] error_io_in_0_a_bits_source;
  wire  error_io_in_0_c_valid;
  wire [2:0] error_io_in_0_c_bits_param;
  wire [3:0] error_io_in_0_c_bits_size;
  wire [4:0] error_io_in_0_c_bits_source;
  wire  error_io_in_0_d_ready;
  wire  error_io_in_0_d_valid;
  wire [2:0] error_io_in_0_d_bits_opcode;
  wire [1:0] error_io_in_0_d_bits_param;
  wire [3:0] error_io_in_0_d_bits_size;
  wire [4:0] error_io_in_0_d_bits_source;
  wire  error_io_in_0_d_bits_sink;
  wire [31:0] error_io_in_0_d_bits_data;
  wire  error_io_in_0_d_bits_error;
  wire  error_TLBuffer_clock;
  wire  error_TLBuffer_reset;
  wire  error_TLBuffer_io_in_0_a_ready;
  wire  error_TLBuffer_io_in_0_a_valid;
  wire [2:0] error_TLBuffer_io_in_0_a_bits_opcode;
  wire [3:0] error_TLBuffer_io_in_0_a_bits_size;
  wire [4:0] error_TLBuffer_io_in_0_a_bits_source;
  wire  error_TLBuffer_io_in_0_d_ready;
  wire  error_TLBuffer_io_in_0_d_valid;
  wire [2:0] error_TLBuffer_io_in_0_d_bits_opcode;
  wire [1:0] error_TLBuffer_io_in_0_d_bits_param;
  wire [3:0] error_TLBuffer_io_in_0_d_bits_size;
  wire [4:0] error_TLBuffer_io_in_0_d_bits_source;
  wire  error_TLBuffer_io_in_0_d_bits_sink;
  wire [31:0] error_TLBuffer_io_in_0_d_bits_data;
  wire  error_TLBuffer_io_in_0_d_bits_error;
  wire  error_TLBuffer_io_out_0_a_ready;
  wire  error_TLBuffer_io_out_0_a_valid;
  wire [2:0] error_TLBuffer_io_out_0_a_bits_opcode;
  wire [3:0] error_TLBuffer_io_out_0_a_bits_size;
  wire [4:0] error_TLBuffer_io_out_0_a_bits_source;
  wire  error_TLBuffer_io_out_0_c_valid;
  wire [2:0] error_TLBuffer_io_out_0_c_bits_param;
  wire [3:0] error_TLBuffer_io_out_0_c_bits_size;
  wire [4:0] error_TLBuffer_io_out_0_c_bits_source;
  wire  error_TLBuffer_io_out_0_d_ready;
  wire  error_TLBuffer_io_out_0_d_valid;
  wire [2:0] error_TLBuffer_io_out_0_d_bits_opcode;
  wire [1:0] error_TLBuffer_io_out_0_d_bits_param;
  wire [3:0] error_TLBuffer_io_out_0_d_bits_size;
  wire [4:0] error_TLBuffer_io_out_0_d_bits_source;
  wire  error_TLBuffer_io_out_0_d_bits_sink;
  wire [31:0] error_TLBuffer_io_out_0_d_bits_data;
  wire  error_TLBuffer_io_out_0_d_bits_error;
  reg [6:0] value;
  reg [31:0] _RAND_0;
  wire  _T_158;
  wire [7:0] _T_160;
  wire [6:0] _T_161;
  wire [6:0] _GEN_0;
  wire  _T_164;
  wire  _T_165;
  IntXbar IntXbar (
    .io_in_0_0(IntXbar_io_in_0_0),
    .io_in_0_1(IntXbar_io_in_0_1),
    .io_out_0_0(IntXbar_io_out_0_0),
    .io_out_0_1(IntXbar_io_out_0_1)
  );
  TLXbar TLXbar (
    .clock(TLXbar_clock),
    .reset(TLXbar_reset),
    .io_in_1_a_ready(TLXbar_io_in_1_a_ready),
    .io_in_1_a_valid(TLXbar_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(TLXbar_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_param(TLXbar_io_in_1_a_bits_param),
    .io_in_1_a_bits_size(TLXbar_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(TLXbar_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(TLXbar_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(TLXbar_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(TLXbar_io_in_1_a_bits_data),
    .io_in_1_d_ready(TLXbar_io_in_1_d_ready),
    .io_in_1_d_valid(TLXbar_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(TLXbar_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_size(TLXbar_io_in_1_d_bits_size),
    .io_in_1_d_bits_source(TLXbar_io_in_1_d_bits_source),
    .io_in_0_a_ready(TLXbar_io_in_0_a_ready),
    .io_in_0_a_valid(TLXbar_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLXbar_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLXbar_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLXbar_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLXbar_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLXbar_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLXbar_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLXbar_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLXbar_io_in_0_d_ready),
    .io_in_0_d_valid(TLXbar_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLXbar_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLXbar_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLXbar_io_in_0_d_bits_source),
    .io_in_0_d_bits_data(TLXbar_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLXbar_io_in_0_d_bits_error),
    .io_out_2_a_ready(TLXbar_io_out_2_a_ready),
    .io_out_2_a_valid(TLXbar_io_out_2_a_valid),
    .io_out_2_a_bits_opcode(TLXbar_io_out_2_a_bits_opcode),
    .io_out_2_a_bits_size(TLXbar_io_out_2_a_bits_size),
    .io_out_2_a_bits_source(TLXbar_io_out_2_a_bits_source),
    .io_out_2_d_ready(TLXbar_io_out_2_d_ready),
    .io_out_2_d_valid(TLXbar_io_out_2_d_valid),
    .io_out_2_d_bits_opcode(TLXbar_io_out_2_d_bits_opcode),
    .io_out_2_d_bits_param(TLXbar_io_out_2_d_bits_param),
    .io_out_2_d_bits_size(TLXbar_io_out_2_d_bits_size),
    .io_out_2_d_bits_source(TLXbar_io_out_2_d_bits_source),
    .io_out_2_d_bits_sink(TLXbar_io_out_2_d_bits_sink),
    .io_out_2_d_bits_data(TLXbar_io_out_2_d_bits_data),
    .io_out_2_d_bits_error(TLXbar_io_out_2_d_bits_error),
    .io_out_1_a_ready(TLXbar_io_out_1_a_ready),
    .io_out_1_a_valid(TLXbar_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLXbar_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(TLXbar_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLXbar_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLXbar_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLXbar_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLXbar_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLXbar_io_out_1_d_ready),
    .io_out_1_d_valid(TLXbar_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLXbar_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(TLXbar_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(TLXbar_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLXbar_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(TLXbar_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(TLXbar_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(TLXbar_io_out_1_d_bits_error),
    .io_out_0_a_ready(TLXbar_io_out_0_a_ready),
    .io_out_0_a_valid(TLXbar_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLXbar_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLXbar_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLXbar_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLXbar_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLXbar_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLXbar_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLXbar_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLXbar_io_out_0_d_ready),
    .io_out_0_d_valid(TLXbar_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLXbar_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLXbar_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLXbar_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLXbar_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLXbar_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLXbar_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLXbar_io_out_0_d_bits_error)
  );
  TLBuffer_1 TLBuffer_1 (
    .clock(TLBuffer_1_clock),
    .reset(TLBuffer_1_reset),
    .io_in_2_a_ready(TLBuffer_1_io_in_2_a_ready),
    .io_in_2_a_valid(TLBuffer_1_io_in_2_a_valid),
    .io_in_2_a_bits_opcode(TLBuffer_1_io_in_2_a_bits_opcode),
    .io_in_2_a_bits_size(TLBuffer_1_io_in_2_a_bits_size),
    .io_in_2_a_bits_source(TLBuffer_1_io_in_2_a_bits_source),
    .io_in_2_d_ready(TLBuffer_1_io_in_2_d_ready),
    .io_in_2_d_valid(TLBuffer_1_io_in_2_d_valid),
    .io_in_2_d_bits_opcode(TLBuffer_1_io_in_2_d_bits_opcode),
    .io_in_2_d_bits_param(TLBuffer_1_io_in_2_d_bits_param),
    .io_in_2_d_bits_size(TLBuffer_1_io_in_2_d_bits_size),
    .io_in_2_d_bits_source(TLBuffer_1_io_in_2_d_bits_source),
    .io_in_2_d_bits_sink(TLBuffer_1_io_in_2_d_bits_sink),
    .io_in_2_d_bits_data(TLBuffer_1_io_in_2_d_bits_data),
    .io_in_2_d_bits_error(TLBuffer_1_io_in_2_d_bits_error),
    .io_in_1_a_ready(TLBuffer_1_io_in_1_a_ready),
    .io_in_1_a_valid(TLBuffer_1_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(TLBuffer_1_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_size(TLBuffer_1_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(TLBuffer_1_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(TLBuffer_1_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(TLBuffer_1_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(TLBuffer_1_io_in_1_a_bits_data),
    .io_in_1_d_ready(TLBuffer_1_io_in_1_d_ready),
    .io_in_1_d_valid(TLBuffer_1_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(TLBuffer_1_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_param(TLBuffer_1_io_in_1_d_bits_param),
    .io_in_1_d_bits_size(TLBuffer_1_io_in_1_d_bits_size),
    .io_in_1_d_bits_source(TLBuffer_1_io_in_1_d_bits_source),
    .io_in_1_d_bits_sink(TLBuffer_1_io_in_1_d_bits_sink),
    .io_in_1_d_bits_data(TLBuffer_1_io_in_1_d_bits_data),
    .io_in_1_d_bits_error(TLBuffer_1_io_in_1_d_bits_error),
    .io_in_0_a_ready(TLBuffer_1_io_in_0_a_ready),
    .io_in_0_a_valid(TLBuffer_1_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLBuffer_1_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLBuffer_1_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLBuffer_1_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLBuffer_1_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLBuffer_1_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLBuffer_1_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLBuffer_1_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLBuffer_1_io_in_0_d_ready),
    .io_in_0_d_valid(TLBuffer_1_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLBuffer_1_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLBuffer_1_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLBuffer_1_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLBuffer_1_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLBuffer_1_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLBuffer_1_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLBuffer_1_io_in_0_d_bits_error),
    .io_out_2_a_ready(TLBuffer_1_io_out_2_a_ready),
    .io_out_2_a_valid(TLBuffer_1_io_out_2_a_valid),
    .io_out_2_a_bits_opcode(TLBuffer_1_io_out_2_a_bits_opcode),
    .io_out_2_a_bits_size(TLBuffer_1_io_out_2_a_bits_size),
    .io_out_2_a_bits_source(TLBuffer_1_io_out_2_a_bits_source),
    .io_out_2_d_ready(TLBuffer_1_io_out_2_d_ready),
    .io_out_2_d_valid(TLBuffer_1_io_out_2_d_valid),
    .io_out_2_d_bits_opcode(TLBuffer_1_io_out_2_d_bits_opcode),
    .io_out_2_d_bits_param(TLBuffer_1_io_out_2_d_bits_param),
    .io_out_2_d_bits_size(TLBuffer_1_io_out_2_d_bits_size),
    .io_out_2_d_bits_source(TLBuffer_1_io_out_2_d_bits_source),
    .io_out_2_d_bits_sink(TLBuffer_1_io_out_2_d_bits_sink),
    .io_out_2_d_bits_data(TLBuffer_1_io_out_2_d_bits_data),
    .io_out_2_d_bits_error(TLBuffer_1_io_out_2_d_bits_error),
    .io_out_1_a_ready(TLBuffer_1_io_out_1_a_ready),
    .io_out_1_a_valid(TLBuffer_1_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLBuffer_1_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(TLBuffer_1_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLBuffer_1_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLBuffer_1_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLBuffer_1_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLBuffer_1_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLBuffer_1_io_out_1_d_ready),
    .io_out_1_d_valid(TLBuffer_1_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLBuffer_1_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(TLBuffer_1_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(TLBuffer_1_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLBuffer_1_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(TLBuffer_1_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(TLBuffer_1_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(TLBuffer_1_io_out_1_d_bits_error),
    .io_out_0_a_ready(TLBuffer_1_io_out_0_a_ready),
    .io_out_0_a_valid(TLBuffer_1_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLBuffer_1_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLBuffer_1_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLBuffer_1_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLBuffer_1_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLBuffer_1_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLBuffer_1_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLBuffer_1_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLBuffer_1_io_out_0_d_ready),
    .io_out_0_d_valid(TLBuffer_1_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLBuffer_1_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLBuffer_1_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLBuffer_1_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLBuffer_1_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLBuffer_1_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLBuffer_1_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLBuffer_1_io_out_0_d_bits_error)
  );
  TLWidthWidget TLWidthWidget (
    .clock(TLWidthWidget_clock),
    .reset(TLWidthWidget_reset),
    .io_in_1_a_ready(TLWidthWidget_io_in_1_a_ready),
    .io_in_1_a_valid(TLWidthWidget_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(TLWidthWidget_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_size(TLWidthWidget_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(TLWidthWidget_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(TLWidthWidget_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(TLWidthWidget_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(TLWidthWidget_io_in_1_a_bits_data),
    .io_in_1_d_ready(TLWidthWidget_io_in_1_d_ready),
    .io_in_1_d_valid(TLWidthWidget_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(TLWidthWidget_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_param(TLWidthWidget_io_in_1_d_bits_param),
    .io_in_1_d_bits_size(TLWidthWidget_io_in_1_d_bits_size),
    .io_in_1_d_bits_source(TLWidthWidget_io_in_1_d_bits_source),
    .io_in_1_d_bits_sink(TLWidthWidget_io_in_1_d_bits_sink),
    .io_in_1_d_bits_data(TLWidthWidget_io_in_1_d_bits_data),
    .io_in_1_d_bits_error(TLWidthWidget_io_in_1_d_bits_error),
    .io_in_0_a_ready(TLWidthWidget_io_in_0_a_ready),
    .io_in_0_a_valid(TLWidthWidget_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLWidthWidget_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLWidthWidget_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLWidthWidget_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLWidthWidget_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLWidthWidget_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLWidthWidget_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLWidthWidget_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLWidthWidget_io_in_0_d_ready),
    .io_in_0_d_valid(TLWidthWidget_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLWidthWidget_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLWidthWidget_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLWidthWidget_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLWidthWidget_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLWidthWidget_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLWidthWidget_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLWidthWidget_io_in_0_d_bits_error),
    .io_out_1_a_ready(TLWidthWidget_io_out_1_a_ready),
    .io_out_1_a_valid(TLWidthWidget_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLWidthWidget_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(TLWidthWidget_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLWidthWidget_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLWidthWidget_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLWidthWidget_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLWidthWidget_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLWidthWidget_io_out_1_d_ready),
    .io_out_1_d_valid(TLWidthWidget_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLWidthWidget_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(TLWidthWidget_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(TLWidthWidget_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLWidthWidget_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(TLWidthWidget_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(TLWidthWidget_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(TLWidthWidget_io_out_1_d_bits_error),
    .io_out_0_a_ready(TLWidthWidget_io_out_0_a_ready),
    .io_out_0_a_valid(TLWidthWidget_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLWidthWidget_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLWidthWidget_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLWidthWidget_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLWidthWidget_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLWidthWidget_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLWidthWidget_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLWidthWidget_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLWidthWidget_io_out_0_d_ready),
    .io_out_0_d_valid(TLWidthWidget_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLWidthWidget_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLWidthWidget_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLWidthWidget_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLWidthWidget_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLWidthWidget_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLWidthWidget_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLWidthWidget_io_out_0_d_bits_error)
  );
  TLSplitter TLSplitter (
    .io_in_1_a_ready(TLSplitter_io_in_1_a_ready),
    .io_in_1_a_valid(TLSplitter_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(TLSplitter_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_param(TLSplitter_io_in_1_a_bits_param),
    .io_in_1_a_bits_size(TLSplitter_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(TLSplitter_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(TLSplitter_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(TLSplitter_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(TLSplitter_io_in_1_a_bits_data),
    .io_in_1_d_ready(TLSplitter_io_in_1_d_ready),
    .io_in_1_d_valid(TLSplitter_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(TLSplitter_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_size(TLSplitter_io_in_1_d_bits_size),
    .io_in_1_d_bits_source(TLSplitter_io_in_1_d_bits_source),
    .io_in_0_a_ready(TLSplitter_io_in_0_a_ready),
    .io_in_0_a_valid(TLSplitter_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLSplitter_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLSplitter_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLSplitter_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLSplitter_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLSplitter_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLSplitter_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLSplitter_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLSplitter_io_in_0_d_ready),
    .io_in_0_d_valid(TLSplitter_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLSplitter_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLSplitter_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLSplitter_io_in_0_d_bits_source),
    .io_in_0_d_bits_data(TLSplitter_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLSplitter_io_in_0_d_bits_error),
    .io_out_1_a_ready(TLSplitter_io_out_1_a_ready),
    .io_out_1_a_valid(TLSplitter_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLSplitter_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_param(TLSplitter_io_out_1_a_bits_param),
    .io_out_1_a_bits_size(TLSplitter_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLSplitter_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLSplitter_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLSplitter_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLSplitter_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLSplitter_io_out_1_d_ready),
    .io_out_1_d_valid(TLSplitter_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLSplitter_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_size(TLSplitter_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLSplitter_io_out_1_d_bits_source),
    .io_out_0_a_ready(TLSplitter_io_out_0_a_ready),
    .io_out_0_a_valid(TLSplitter_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLSplitter_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLSplitter_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLSplitter_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLSplitter_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLSplitter_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLSplitter_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLSplitter_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLSplitter_io_out_0_d_ready),
    .io_out_0_d_valid(TLSplitter_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLSplitter_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(TLSplitter_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLSplitter_io_out_0_d_bits_source),
    .io_out_0_d_bits_data(TLSplitter_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLSplitter_io_out_0_d_bits_error)
  );
  TLFIFOFixer TLFIFOFixer (
    .io_in_0_a_ready(TLFIFOFixer_io_in_0_a_ready),
    .io_in_0_a_valid(TLFIFOFixer_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLFIFOFixer_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLFIFOFixer_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLFIFOFixer_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLFIFOFixer_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLFIFOFixer_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLFIFOFixer_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLFIFOFixer_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLFIFOFixer_io_in_0_d_ready),
    .io_in_0_d_valid(TLFIFOFixer_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLFIFOFixer_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLFIFOFixer_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLFIFOFixer_io_in_0_d_bits_source),
    .io_in_0_d_bits_data(TLFIFOFixer_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLFIFOFixer_io_in_0_d_bits_error),
    .io_out_0_a_ready(TLFIFOFixer_io_out_0_a_ready),
    .io_out_0_a_valid(TLFIFOFixer_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLFIFOFixer_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLFIFOFixer_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLFIFOFixer_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLFIFOFixer_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLFIFOFixer_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLFIFOFixer_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLFIFOFixer_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLFIFOFixer_io_out_0_d_ready),
    .io_out_0_d_valid(TLFIFOFixer_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLFIFOFixer_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(TLFIFOFixer_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLFIFOFixer_io_out_0_d_bits_source),
    .io_out_0_d_bits_data(TLFIFOFixer_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLFIFOFixer_io_out_0_d_bits_error)
  );
  TLFIFOFixer_1 TLFIFOFixer_1 (
    .clock(TLFIFOFixer_1_clock),
    .reset(TLFIFOFixer_1_reset),
    .io_in_0_a_ready(TLFIFOFixer_1_io_in_0_a_ready),
    .io_in_0_a_valid(TLFIFOFixer_1_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLFIFOFixer_1_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLFIFOFixer_1_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLFIFOFixer_1_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLFIFOFixer_1_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLFIFOFixer_1_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLFIFOFixer_1_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLFIFOFixer_1_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLFIFOFixer_1_io_in_0_d_ready),
    .io_in_0_d_valid(TLFIFOFixer_1_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLFIFOFixer_1_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLFIFOFixer_1_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLFIFOFixer_1_io_in_0_d_bits_source),
    .io_out_0_a_ready(TLFIFOFixer_1_io_out_0_a_ready),
    .io_out_0_a_valid(TLFIFOFixer_1_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLFIFOFixer_1_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLFIFOFixer_1_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLFIFOFixer_1_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLFIFOFixer_1_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLFIFOFixer_1_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLFIFOFixer_1_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLFIFOFixer_1_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLFIFOFixer_1_io_out_0_d_ready),
    .io_out_0_d_valid(TLFIFOFixer_1_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLFIFOFixer_1_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(TLFIFOFixer_1_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLFIFOFixer_1_io_out_0_d_bits_source)
  );
  TLXbar_1 TLXbar_1 (
    .clock(TLXbar_1_clock),
    .reset(TLXbar_1_reset),
    .io_in_0_a_ready(TLXbar_1_io_in_0_a_ready),
    .io_in_0_a_valid(TLXbar_1_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLXbar_1_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLXbar_1_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLXbar_1_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLXbar_1_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLXbar_1_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLXbar_1_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLXbar_1_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLXbar_1_io_in_0_d_ready),
    .io_in_0_d_valid(TLXbar_1_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLXbar_1_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLXbar_1_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLXbar_1_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLXbar_1_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLXbar_1_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLXbar_1_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLXbar_1_io_in_0_d_bits_error),
    .io_out_4_a_ready(TLXbar_1_io_out_4_a_ready),
    .io_out_4_a_valid(TLXbar_1_io_out_4_a_valid),
    .io_out_4_a_bits_opcode(TLXbar_1_io_out_4_a_bits_opcode),
    .io_out_4_a_bits_param(TLXbar_1_io_out_4_a_bits_param),
    .io_out_4_a_bits_size(TLXbar_1_io_out_4_a_bits_size),
    .io_out_4_a_bits_source(TLXbar_1_io_out_4_a_bits_source),
    .io_out_4_a_bits_address(TLXbar_1_io_out_4_a_bits_address),
    .io_out_4_a_bits_mask(TLXbar_1_io_out_4_a_bits_mask),
    .io_out_4_a_bits_data(TLXbar_1_io_out_4_a_bits_data),
    .io_out_4_d_ready(TLXbar_1_io_out_4_d_ready),
    .io_out_4_d_valid(TLXbar_1_io_out_4_d_valid),
    .io_out_4_d_bits_opcode(TLXbar_1_io_out_4_d_bits_opcode),
    .io_out_4_d_bits_param(TLXbar_1_io_out_4_d_bits_param),
    .io_out_4_d_bits_size(TLXbar_1_io_out_4_d_bits_size),
    .io_out_4_d_bits_source(TLXbar_1_io_out_4_d_bits_source),
    .io_out_4_d_bits_sink(TLXbar_1_io_out_4_d_bits_sink),
    .io_out_4_d_bits_data(TLXbar_1_io_out_4_d_bits_data),
    .io_out_4_d_bits_error(TLXbar_1_io_out_4_d_bits_error),
    .io_out_3_a_ready(TLXbar_1_io_out_3_a_ready),
    .io_out_3_a_valid(TLXbar_1_io_out_3_a_valid),
    .io_out_3_a_bits_opcode(TLXbar_1_io_out_3_a_bits_opcode),
    .io_out_3_a_bits_size(TLXbar_1_io_out_3_a_bits_size),
    .io_out_3_a_bits_source(TLXbar_1_io_out_3_a_bits_source),
    .io_out_3_a_bits_address(TLXbar_1_io_out_3_a_bits_address),
    .io_out_3_a_bits_mask(TLXbar_1_io_out_3_a_bits_mask),
    .io_out_3_d_ready(TLXbar_1_io_out_3_d_ready),
    .io_out_3_d_valid(TLXbar_1_io_out_3_d_valid),
    .io_out_3_d_bits_opcode(TLXbar_1_io_out_3_d_bits_opcode),
    .io_out_3_d_bits_param(TLXbar_1_io_out_3_d_bits_param),
    .io_out_3_d_bits_size(TLXbar_1_io_out_3_d_bits_size),
    .io_out_3_d_bits_source(TLXbar_1_io_out_3_d_bits_source),
    .io_out_3_d_bits_sink(TLXbar_1_io_out_3_d_bits_sink),
    .io_out_3_d_bits_data(TLXbar_1_io_out_3_d_bits_data),
    .io_out_3_d_bits_error(TLXbar_1_io_out_3_d_bits_error),
    .io_out_2_a_ready(TLXbar_1_io_out_2_a_ready),
    .io_out_2_a_valid(TLXbar_1_io_out_2_a_valid),
    .io_out_2_a_bits_opcode(TLXbar_1_io_out_2_a_bits_opcode),
    .io_out_2_a_bits_size(TLXbar_1_io_out_2_a_bits_size),
    .io_out_2_a_bits_source(TLXbar_1_io_out_2_a_bits_source),
    .io_out_2_a_bits_address(TLXbar_1_io_out_2_a_bits_address),
    .io_out_2_a_bits_mask(TLXbar_1_io_out_2_a_bits_mask),
    .io_out_2_a_bits_data(TLXbar_1_io_out_2_a_bits_data),
    .io_out_2_d_ready(TLXbar_1_io_out_2_d_ready),
    .io_out_2_d_valid(TLXbar_1_io_out_2_d_valid),
    .io_out_2_d_bits_opcode(TLXbar_1_io_out_2_d_bits_opcode),
    .io_out_2_d_bits_param(TLXbar_1_io_out_2_d_bits_param),
    .io_out_2_d_bits_size(TLXbar_1_io_out_2_d_bits_size),
    .io_out_2_d_bits_source(TLXbar_1_io_out_2_d_bits_source),
    .io_out_2_d_bits_sink(TLXbar_1_io_out_2_d_bits_sink),
    .io_out_2_d_bits_data(TLXbar_1_io_out_2_d_bits_data),
    .io_out_2_d_bits_error(TLXbar_1_io_out_2_d_bits_error),
    .io_out_1_a_ready(TLXbar_1_io_out_1_a_ready),
    .io_out_1_a_valid(TLXbar_1_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLXbar_1_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(TLXbar_1_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLXbar_1_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLXbar_1_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLXbar_1_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLXbar_1_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLXbar_1_io_out_1_d_ready),
    .io_out_1_d_valid(TLXbar_1_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLXbar_1_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(TLXbar_1_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(TLXbar_1_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLXbar_1_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(TLXbar_1_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(TLXbar_1_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(TLXbar_1_io_out_1_d_bits_error),
    .io_out_0_a_ready(TLXbar_1_io_out_0_a_ready),
    .io_out_0_a_valid(TLXbar_1_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLXbar_1_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(TLXbar_1_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLXbar_1_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLXbar_1_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLXbar_1_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLXbar_1_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLXbar_1_io_out_0_d_ready),
    .io_out_0_d_valid(TLXbar_1_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLXbar_1_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLXbar_1_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLXbar_1_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLXbar_1_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLXbar_1_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLXbar_1_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLXbar_1_io_out_0_d_bits_error)
  );
  TLBuffer_2 TLBuffer_2 (
    .clock(TLBuffer_2_clock),
    .reset(TLBuffer_2_reset),
    .io_in_0_a_ready(TLBuffer_2_io_in_0_a_ready),
    .io_in_0_a_valid(TLBuffer_2_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLBuffer_2_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLBuffer_2_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLBuffer_2_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLBuffer_2_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLBuffer_2_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLBuffer_2_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLBuffer_2_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLBuffer_2_io_in_0_d_ready),
    .io_in_0_d_valid(TLBuffer_2_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLBuffer_2_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLBuffer_2_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLBuffer_2_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLBuffer_2_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLBuffer_2_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLBuffer_2_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLBuffer_2_io_in_0_d_bits_error),
    .io_out_0_a_ready(TLBuffer_2_io_out_0_a_ready),
    .io_out_0_a_valid(TLBuffer_2_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLBuffer_2_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLBuffer_2_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLBuffer_2_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLBuffer_2_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLBuffer_2_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLBuffer_2_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLBuffer_2_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLBuffer_2_io_out_0_d_ready),
    .io_out_0_d_valid(TLBuffer_2_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLBuffer_2_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLBuffer_2_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLBuffer_2_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLBuffer_2_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLBuffer_2_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLBuffer_2_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLBuffer_2_io_out_0_d_bits_error)
  );
  TLBuffer_3 TLBuffer_3 (
    .io_in_4_a_ready(TLBuffer_3_io_in_4_a_ready),
    .io_in_4_a_valid(TLBuffer_3_io_in_4_a_valid),
    .io_in_4_a_bits_opcode(TLBuffer_3_io_in_4_a_bits_opcode),
    .io_in_4_a_bits_param(TLBuffer_3_io_in_4_a_bits_param),
    .io_in_4_a_bits_size(TLBuffer_3_io_in_4_a_bits_size),
    .io_in_4_a_bits_source(TLBuffer_3_io_in_4_a_bits_source),
    .io_in_4_a_bits_address(TLBuffer_3_io_in_4_a_bits_address),
    .io_in_4_a_bits_mask(TLBuffer_3_io_in_4_a_bits_mask),
    .io_in_4_a_bits_data(TLBuffer_3_io_in_4_a_bits_data),
    .io_in_4_d_ready(TLBuffer_3_io_in_4_d_ready),
    .io_in_4_d_valid(TLBuffer_3_io_in_4_d_valid),
    .io_in_4_d_bits_opcode(TLBuffer_3_io_in_4_d_bits_opcode),
    .io_in_4_d_bits_param(TLBuffer_3_io_in_4_d_bits_param),
    .io_in_4_d_bits_size(TLBuffer_3_io_in_4_d_bits_size),
    .io_in_4_d_bits_source(TLBuffer_3_io_in_4_d_bits_source),
    .io_in_4_d_bits_sink(TLBuffer_3_io_in_4_d_bits_sink),
    .io_in_4_d_bits_data(TLBuffer_3_io_in_4_d_bits_data),
    .io_in_4_d_bits_error(TLBuffer_3_io_in_4_d_bits_error),
    .io_in_3_a_ready(TLBuffer_3_io_in_3_a_ready),
    .io_in_3_a_valid(TLBuffer_3_io_in_3_a_valid),
    .io_in_3_a_bits_opcode(TLBuffer_3_io_in_3_a_bits_opcode),
    .io_in_3_a_bits_size(TLBuffer_3_io_in_3_a_bits_size),
    .io_in_3_a_bits_source(TLBuffer_3_io_in_3_a_bits_source),
    .io_in_3_a_bits_address(TLBuffer_3_io_in_3_a_bits_address),
    .io_in_3_a_bits_mask(TLBuffer_3_io_in_3_a_bits_mask),
    .io_in_3_d_ready(TLBuffer_3_io_in_3_d_ready),
    .io_in_3_d_valid(TLBuffer_3_io_in_3_d_valid),
    .io_in_3_d_bits_opcode(TLBuffer_3_io_in_3_d_bits_opcode),
    .io_in_3_d_bits_param(TLBuffer_3_io_in_3_d_bits_param),
    .io_in_3_d_bits_size(TLBuffer_3_io_in_3_d_bits_size),
    .io_in_3_d_bits_source(TLBuffer_3_io_in_3_d_bits_source),
    .io_in_3_d_bits_sink(TLBuffer_3_io_in_3_d_bits_sink),
    .io_in_3_d_bits_data(TLBuffer_3_io_in_3_d_bits_data),
    .io_in_3_d_bits_error(TLBuffer_3_io_in_3_d_bits_error),
    .io_in_2_a_ready(TLBuffer_3_io_in_2_a_ready),
    .io_in_2_a_valid(TLBuffer_3_io_in_2_a_valid),
    .io_in_2_a_bits_opcode(TLBuffer_3_io_in_2_a_bits_opcode),
    .io_in_2_a_bits_size(TLBuffer_3_io_in_2_a_bits_size),
    .io_in_2_a_bits_source(TLBuffer_3_io_in_2_a_bits_source),
    .io_in_2_a_bits_address(TLBuffer_3_io_in_2_a_bits_address),
    .io_in_2_a_bits_mask(TLBuffer_3_io_in_2_a_bits_mask),
    .io_in_2_a_bits_data(TLBuffer_3_io_in_2_a_bits_data),
    .io_in_2_d_ready(TLBuffer_3_io_in_2_d_ready),
    .io_in_2_d_valid(TLBuffer_3_io_in_2_d_valid),
    .io_in_2_d_bits_opcode(TLBuffer_3_io_in_2_d_bits_opcode),
    .io_in_2_d_bits_param(TLBuffer_3_io_in_2_d_bits_param),
    .io_in_2_d_bits_size(TLBuffer_3_io_in_2_d_bits_size),
    .io_in_2_d_bits_source(TLBuffer_3_io_in_2_d_bits_source),
    .io_in_2_d_bits_sink(TLBuffer_3_io_in_2_d_bits_sink),
    .io_in_2_d_bits_data(TLBuffer_3_io_in_2_d_bits_data),
    .io_in_2_d_bits_error(TLBuffer_3_io_in_2_d_bits_error),
    .io_in_1_a_ready(TLBuffer_3_io_in_1_a_ready),
    .io_in_1_a_valid(TLBuffer_3_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(TLBuffer_3_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_size(TLBuffer_3_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(TLBuffer_3_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(TLBuffer_3_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(TLBuffer_3_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(TLBuffer_3_io_in_1_a_bits_data),
    .io_in_1_d_ready(TLBuffer_3_io_in_1_d_ready),
    .io_in_1_d_valid(TLBuffer_3_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(TLBuffer_3_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_param(TLBuffer_3_io_in_1_d_bits_param),
    .io_in_1_d_bits_size(TLBuffer_3_io_in_1_d_bits_size),
    .io_in_1_d_bits_source(TLBuffer_3_io_in_1_d_bits_source),
    .io_in_1_d_bits_sink(TLBuffer_3_io_in_1_d_bits_sink),
    .io_in_1_d_bits_data(TLBuffer_3_io_in_1_d_bits_data),
    .io_in_1_d_bits_error(TLBuffer_3_io_in_1_d_bits_error),
    .io_in_0_a_ready(TLBuffer_3_io_in_0_a_ready),
    .io_in_0_a_valid(TLBuffer_3_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLBuffer_3_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(TLBuffer_3_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLBuffer_3_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLBuffer_3_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLBuffer_3_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLBuffer_3_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLBuffer_3_io_in_0_d_ready),
    .io_in_0_d_valid(TLBuffer_3_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLBuffer_3_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLBuffer_3_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLBuffer_3_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLBuffer_3_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLBuffer_3_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLBuffer_3_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLBuffer_3_io_in_0_d_bits_error),
    .io_out_4_a_ready(TLBuffer_3_io_out_4_a_ready),
    .io_out_4_a_valid(TLBuffer_3_io_out_4_a_valid),
    .io_out_4_a_bits_opcode(TLBuffer_3_io_out_4_a_bits_opcode),
    .io_out_4_a_bits_param(TLBuffer_3_io_out_4_a_bits_param),
    .io_out_4_a_bits_size(TLBuffer_3_io_out_4_a_bits_size),
    .io_out_4_a_bits_source(TLBuffer_3_io_out_4_a_bits_source),
    .io_out_4_a_bits_address(TLBuffer_3_io_out_4_a_bits_address),
    .io_out_4_a_bits_mask(TLBuffer_3_io_out_4_a_bits_mask),
    .io_out_4_a_bits_data(TLBuffer_3_io_out_4_a_bits_data),
    .io_out_4_d_ready(TLBuffer_3_io_out_4_d_ready),
    .io_out_4_d_valid(TLBuffer_3_io_out_4_d_valid),
    .io_out_4_d_bits_opcode(TLBuffer_3_io_out_4_d_bits_opcode),
    .io_out_4_d_bits_param(TLBuffer_3_io_out_4_d_bits_param),
    .io_out_4_d_bits_size(TLBuffer_3_io_out_4_d_bits_size),
    .io_out_4_d_bits_source(TLBuffer_3_io_out_4_d_bits_source),
    .io_out_4_d_bits_sink(TLBuffer_3_io_out_4_d_bits_sink),
    .io_out_4_d_bits_data(TLBuffer_3_io_out_4_d_bits_data),
    .io_out_4_d_bits_error(TLBuffer_3_io_out_4_d_bits_error),
    .io_out_3_a_ready(TLBuffer_3_io_out_3_a_ready),
    .io_out_3_a_valid(TLBuffer_3_io_out_3_a_valid),
    .io_out_3_a_bits_opcode(TLBuffer_3_io_out_3_a_bits_opcode),
    .io_out_3_a_bits_size(TLBuffer_3_io_out_3_a_bits_size),
    .io_out_3_a_bits_source(TLBuffer_3_io_out_3_a_bits_source),
    .io_out_3_a_bits_address(TLBuffer_3_io_out_3_a_bits_address),
    .io_out_3_a_bits_mask(TLBuffer_3_io_out_3_a_bits_mask),
    .io_out_3_d_ready(TLBuffer_3_io_out_3_d_ready),
    .io_out_3_d_valid(TLBuffer_3_io_out_3_d_valid),
    .io_out_3_d_bits_opcode(TLBuffer_3_io_out_3_d_bits_opcode),
    .io_out_3_d_bits_param(TLBuffer_3_io_out_3_d_bits_param),
    .io_out_3_d_bits_size(TLBuffer_3_io_out_3_d_bits_size),
    .io_out_3_d_bits_source(TLBuffer_3_io_out_3_d_bits_source),
    .io_out_3_d_bits_sink(TLBuffer_3_io_out_3_d_bits_sink),
    .io_out_3_d_bits_data(TLBuffer_3_io_out_3_d_bits_data),
    .io_out_3_d_bits_error(TLBuffer_3_io_out_3_d_bits_error),
    .io_out_2_a_ready(TLBuffer_3_io_out_2_a_ready),
    .io_out_2_a_valid(TLBuffer_3_io_out_2_a_valid),
    .io_out_2_a_bits_opcode(TLBuffer_3_io_out_2_a_bits_opcode),
    .io_out_2_a_bits_size(TLBuffer_3_io_out_2_a_bits_size),
    .io_out_2_a_bits_source(TLBuffer_3_io_out_2_a_bits_source),
    .io_out_2_a_bits_address(TLBuffer_3_io_out_2_a_bits_address),
    .io_out_2_a_bits_mask(TLBuffer_3_io_out_2_a_bits_mask),
    .io_out_2_a_bits_data(TLBuffer_3_io_out_2_a_bits_data),
    .io_out_2_d_ready(TLBuffer_3_io_out_2_d_ready),
    .io_out_2_d_valid(TLBuffer_3_io_out_2_d_valid),
    .io_out_2_d_bits_opcode(TLBuffer_3_io_out_2_d_bits_opcode),
    .io_out_2_d_bits_param(TLBuffer_3_io_out_2_d_bits_param),
    .io_out_2_d_bits_size(TLBuffer_3_io_out_2_d_bits_size),
    .io_out_2_d_bits_source(TLBuffer_3_io_out_2_d_bits_source),
    .io_out_2_d_bits_sink(TLBuffer_3_io_out_2_d_bits_sink),
    .io_out_2_d_bits_data(TLBuffer_3_io_out_2_d_bits_data),
    .io_out_2_d_bits_error(TLBuffer_3_io_out_2_d_bits_error),
    .io_out_1_a_ready(TLBuffer_3_io_out_1_a_ready),
    .io_out_1_a_valid(TLBuffer_3_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLBuffer_3_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(TLBuffer_3_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLBuffer_3_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLBuffer_3_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLBuffer_3_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLBuffer_3_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLBuffer_3_io_out_1_d_ready),
    .io_out_1_d_valid(TLBuffer_3_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLBuffer_3_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(TLBuffer_3_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(TLBuffer_3_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLBuffer_3_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(TLBuffer_3_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(TLBuffer_3_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(TLBuffer_3_io_out_1_d_bits_error),
    .io_out_0_a_ready(TLBuffer_3_io_out_0_a_ready),
    .io_out_0_a_valid(TLBuffer_3_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLBuffer_3_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(TLBuffer_3_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLBuffer_3_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLBuffer_3_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLBuffer_3_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLBuffer_3_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLBuffer_3_io_out_0_d_ready),
    .io_out_0_d_valid(TLBuffer_3_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLBuffer_3_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLBuffer_3_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLBuffer_3_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLBuffer_3_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLBuffer_3_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLBuffer_3_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLBuffer_3_io_out_0_d_bits_error)
  );
  TLFragmenter_1 TLFragmenter_1 (
    .clock(TLFragmenter_1_clock),
    .reset(TLFragmenter_1_reset),
    .io_in_3_a_ready(TLFragmenter_1_io_in_3_a_ready),
    .io_in_3_a_valid(TLFragmenter_1_io_in_3_a_valid),
    .io_in_3_a_bits_opcode(TLFragmenter_1_io_in_3_a_bits_opcode),
    .io_in_3_a_bits_size(TLFragmenter_1_io_in_3_a_bits_size),
    .io_in_3_a_bits_source(TLFragmenter_1_io_in_3_a_bits_source),
    .io_in_3_a_bits_address(TLFragmenter_1_io_in_3_a_bits_address),
    .io_in_3_a_bits_mask(TLFragmenter_1_io_in_3_a_bits_mask),
    .io_in_3_d_ready(TLFragmenter_1_io_in_3_d_ready),
    .io_in_3_d_valid(TLFragmenter_1_io_in_3_d_valid),
    .io_in_3_d_bits_opcode(TLFragmenter_1_io_in_3_d_bits_opcode),
    .io_in_3_d_bits_param(TLFragmenter_1_io_in_3_d_bits_param),
    .io_in_3_d_bits_size(TLFragmenter_1_io_in_3_d_bits_size),
    .io_in_3_d_bits_source(TLFragmenter_1_io_in_3_d_bits_source),
    .io_in_3_d_bits_sink(TLFragmenter_1_io_in_3_d_bits_sink),
    .io_in_3_d_bits_data(TLFragmenter_1_io_in_3_d_bits_data),
    .io_in_3_d_bits_error(TLFragmenter_1_io_in_3_d_bits_error),
    .io_in_2_a_ready(TLFragmenter_1_io_in_2_a_ready),
    .io_in_2_a_valid(TLFragmenter_1_io_in_2_a_valid),
    .io_in_2_a_bits_opcode(TLFragmenter_1_io_in_2_a_bits_opcode),
    .io_in_2_a_bits_size(TLFragmenter_1_io_in_2_a_bits_size),
    .io_in_2_a_bits_source(TLFragmenter_1_io_in_2_a_bits_source),
    .io_in_2_a_bits_address(TLFragmenter_1_io_in_2_a_bits_address),
    .io_in_2_a_bits_mask(TLFragmenter_1_io_in_2_a_bits_mask),
    .io_in_2_a_bits_data(TLFragmenter_1_io_in_2_a_bits_data),
    .io_in_2_d_ready(TLFragmenter_1_io_in_2_d_ready),
    .io_in_2_d_valid(TLFragmenter_1_io_in_2_d_valid),
    .io_in_2_d_bits_opcode(TLFragmenter_1_io_in_2_d_bits_opcode),
    .io_in_2_d_bits_param(TLFragmenter_1_io_in_2_d_bits_param),
    .io_in_2_d_bits_size(TLFragmenter_1_io_in_2_d_bits_size),
    .io_in_2_d_bits_source(TLFragmenter_1_io_in_2_d_bits_source),
    .io_in_2_d_bits_sink(TLFragmenter_1_io_in_2_d_bits_sink),
    .io_in_2_d_bits_data(TLFragmenter_1_io_in_2_d_bits_data),
    .io_in_2_d_bits_error(TLFragmenter_1_io_in_2_d_bits_error),
    .io_in_1_a_ready(TLFragmenter_1_io_in_1_a_ready),
    .io_in_1_a_valid(TLFragmenter_1_io_in_1_a_valid),
    .io_in_1_a_bits_opcode(TLFragmenter_1_io_in_1_a_bits_opcode),
    .io_in_1_a_bits_size(TLFragmenter_1_io_in_1_a_bits_size),
    .io_in_1_a_bits_source(TLFragmenter_1_io_in_1_a_bits_source),
    .io_in_1_a_bits_address(TLFragmenter_1_io_in_1_a_bits_address),
    .io_in_1_a_bits_mask(TLFragmenter_1_io_in_1_a_bits_mask),
    .io_in_1_a_bits_data(TLFragmenter_1_io_in_1_a_bits_data),
    .io_in_1_d_ready(TLFragmenter_1_io_in_1_d_ready),
    .io_in_1_d_valid(TLFragmenter_1_io_in_1_d_valid),
    .io_in_1_d_bits_opcode(TLFragmenter_1_io_in_1_d_bits_opcode),
    .io_in_1_d_bits_param(TLFragmenter_1_io_in_1_d_bits_param),
    .io_in_1_d_bits_size(TLFragmenter_1_io_in_1_d_bits_size),
    .io_in_1_d_bits_source(TLFragmenter_1_io_in_1_d_bits_source),
    .io_in_1_d_bits_sink(TLFragmenter_1_io_in_1_d_bits_sink),
    .io_in_1_d_bits_data(TLFragmenter_1_io_in_1_d_bits_data),
    .io_in_1_d_bits_error(TLFragmenter_1_io_in_1_d_bits_error),
    .io_in_0_a_ready(TLFragmenter_1_io_in_0_a_ready),
    .io_in_0_a_valid(TLFragmenter_1_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLFragmenter_1_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(TLFragmenter_1_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLFragmenter_1_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLFragmenter_1_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLFragmenter_1_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLFragmenter_1_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLFragmenter_1_io_in_0_d_ready),
    .io_in_0_d_valid(TLFragmenter_1_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLFragmenter_1_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLFragmenter_1_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLFragmenter_1_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLFragmenter_1_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLFragmenter_1_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLFragmenter_1_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLFragmenter_1_io_in_0_d_bits_error),
    .io_out_3_a_ready(TLFragmenter_1_io_out_3_a_ready),
    .io_out_3_a_valid(TLFragmenter_1_io_out_3_a_valid),
    .io_out_3_a_bits_size(TLFragmenter_1_io_out_3_a_bits_size),
    .io_out_3_a_bits_source(TLFragmenter_1_io_out_3_a_bits_source),
    .io_out_3_a_bits_address(TLFragmenter_1_io_out_3_a_bits_address),
    .io_out_3_d_ready(TLFragmenter_1_io_out_3_d_ready),
    .io_out_3_d_valid(TLFragmenter_1_io_out_3_d_valid),
    .io_out_3_d_bits_opcode(TLFragmenter_1_io_out_3_d_bits_opcode),
    .io_out_3_d_bits_param(TLFragmenter_1_io_out_3_d_bits_param),
    .io_out_3_d_bits_size(TLFragmenter_1_io_out_3_d_bits_size),
    .io_out_3_d_bits_source(TLFragmenter_1_io_out_3_d_bits_source),
    .io_out_3_d_bits_sink(TLFragmenter_1_io_out_3_d_bits_sink),
    .io_out_3_d_bits_data(TLFragmenter_1_io_out_3_d_bits_data),
    .io_out_3_d_bits_error(TLFragmenter_1_io_out_3_d_bits_error),
    .io_out_2_a_ready(TLFragmenter_1_io_out_2_a_ready),
    .io_out_2_a_valid(TLFragmenter_1_io_out_2_a_valid),
    .io_out_2_a_bits_opcode(TLFragmenter_1_io_out_2_a_bits_opcode),
    .io_out_2_a_bits_size(TLFragmenter_1_io_out_2_a_bits_size),
    .io_out_2_a_bits_source(TLFragmenter_1_io_out_2_a_bits_source),
    .io_out_2_a_bits_address(TLFragmenter_1_io_out_2_a_bits_address),
    .io_out_2_a_bits_mask(TLFragmenter_1_io_out_2_a_bits_mask),
    .io_out_2_a_bits_data(TLFragmenter_1_io_out_2_a_bits_data),
    .io_out_2_d_ready(TLFragmenter_1_io_out_2_d_ready),
    .io_out_2_d_valid(TLFragmenter_1_io_out_2_d_valid),
    .io_out_2_d_bits_opcode(TLFragmenter_1_io_out_2_d_bits_opcode),
    .io_out_2_d_bits_param(TLFragmenter_1_io_out_2_d_bits_param),
    .io_out_2_d_bits_size(TLFragmenter_1_io_out_2_d_bits_size),
    .io_out_2_d_bits_source(TLFragmenter_1_io_out_2_d_bits_source),
    .io_out_2_d_bits_sink(TLFragmenter_1_io_out_2_d_bits_sink),
    .io_out_2_d_bits_data(TLFragmenter_1_io_out_2_d_bits_data),
    .io_out_2_d_bits_error(TLFragmenter_1_io_out_2_d_bits_error),
    .io_out_1_a_ready(TLFragmenter_1_io_out_1_a_ready),
    .io_out_1_a_valid(TLFragmenter_1_io_out_1_a_valid),
    .io_out_1_a_bits_opcode(TLFragmenter_1_io_out_1_a_bits_opcode),
    .io_out_1_a_bits_size(TLFragmenter_1_io_out_1_a_bits_size),
    .io_out_1_a_bits_source(TLFragmenter_1_io_out_1_a_bits_source),
    .io_out_1_a_bits_address(TLFragmenter_1_io_out_1_a_bits_address),
    .io_out_1_a_bits_mask(TLFragmenter_1_io_out_1_a_bits_mask),
    .io_out_1_a_bits_data(TLFragmenter_1_io_out_1_a_bits_data),
    .io_out_1_d_ready(TLFragmenter_1_io_out_1_d_ready),
    .io_out_1_d_valid(TLFragmenter_1_io_out_1_d_valid),
    .io_out_1_d_bits_opcode(TLFragmenter_1_io_out_1_d_bits_opcode),
    .io_out_1_d_bits_param(TLFragmenter_1_io_out_1_d_bits_param),
    .io_out_1_d_bits_size(TLFragmenter_1_io_out_1_d_bits_size),
    .io_out_1_d_bits_source(TLFragmenter_1_io_out_1_d_bits_source),
    .io_out_1_d_bits_sink(TLFragmenter_1_io_out_1_d_bits_sink),
    .io_out_1_d_bits_data(TLFragmenter_1_io_out_1_d_bits_data),
    .io_out_1_d_bits_error(TLFragmenter_1_io_out_1_d_bits_error),
    .io_out_0_a_ready(TLFragmenter_1_io_out_0_a_ready),
    .io_out_0_a_valid(TLFragmenter_1_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLFragmenter_1_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(TLFragmenter_1_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLFragmenter_1_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLFragmenter_1_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLFragmenter_1_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLFragmenter_1_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLFragmenter_1_io_out_0_d_ready),
    .io_out_0_d_valid(TLFragmenter_1_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLFragmenter_1_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLFragmenter_1_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLFragmenter_1_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLFragmenter_1_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLFragmenter_1_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLFragmenter_1_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLFragmenter_1_io_out_0_d_bits_error)
  );
  TLAtomicAutomata TLAtomicAutomata (
    .clock(TLAtomicAutomata_clock),
    .reset(TLAtomicAutomata_reset),
    .io_in_0_a_ready(TLAtomicAutomata_io_in_0_a_ready),
    .io_in_0_a_valid(TLAtomicAutomata_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLAtomicAutomata_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLAtomicAutomata_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLAtomicAutomata_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLAtomicAutomata_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLAtomicAutomata_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLAtomicAutomata_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLAtomicAutomata_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLAtomicAutomata_io_in_0_d_ready),
    .io_in_0_d_valid(TLAtomicAutomata_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLAtomicAutomata_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLAtomicAutomata_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLAtomicAutomata_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLAtomicAutomata_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLAtomicAutomata_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLAtomicAutomata_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLAtomicAutomata_io_in_0_d_bits_error),
    .io_out_0_a_ready(TLAtomicAutomata_io_out_0_a_ready),
    .io_out_0_a_valid(TLAtomicAutomata_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLAtomicAutomata_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLAtomicAutomata_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLAtomicAutomata_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLAtomicAutomata_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLAtomicAutomata_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLAtomicAutomata_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLAtomicAutomata_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLAtomicAutomata_io_out_0_d_ready),
    .io_out_0_d_valid(TLAtomicAutomata_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLAtomicAutomata_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(TLAtomicAutomata_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(TLAtomicAutomata_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLAtomicAutomata_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(TLAtomicAutomata_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(TLAtomicAutomata_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLAtomicAutomata_io_out_0_d_bits_error)
  );
  TLPLIC_plic plic (
    .clock(plic_clock),
    .reset(plic_reset),
    .io_tl_in_0_a_ready(plic_io_tl_in_0_a_ready),
    .io_tl_in_0_a_valid(plic_io_tl_in_0_a_valid),
    .io_tl_in_0_a_bits_opcode(plic_io_tl_in_0_a_bits_opcode),
    .io_tl_in_0_a_bits_size(plic_io_tl_in_0_a_bits_size),
    .io_tl_in_0_a_bits_source(plic_io_tl_in_0_a_bits_source),
    .io_tl_in_0_a_bits_address(plic_io_tl_in_0_a_bits_address),
    .io_tl_in_0_a_bits_mask(plic_io_tl_in_0_a_bits_mask),
    .io_tl_in_0_a_bits_data(plic_io_tl_in_0_a_bits_data),
    .io_tl_in_0_d_ready(plic_io_tl_in_0_d_ready),
    .io_tl_in_0_d_valid(plic_io_tl_in_0_d_valid),
    .io_tl_in_0_d_bits_opcode(plic_io_tl_in_0_d_bits_opcode),
    .io_tl_in_0_d_bits_param(plic_io_tl_in_0_d_bits_param),
    .io_tl_in_0_d_bits_size(plic_io_tl_in_0_d_bits_size),
    .io_tl_in_0_d_bits_source(plic_io_tl_in_0_d_bits_source),
    .io_tl_in_0_d_bits_sink(plic_io_tl_in_0_d_bits_sink),
    .io_tl_in_0_d_bits_data(plic_io_tl_in_0_d_bits_data),
    .io_tl_in_0_d_bits_error(plic_io_tl_in_0_d_bits_error),
    .io_devices_0_0(plic_io_devices_0_0),
    .io_devices_0_1(plic_io_devices_0_1),
    .io_harts_0_0(plic_io_harts_0_0)
  );
  CoreplexLocalInterrupter_clint clint (
    .clock(clint_clock),
    .reset(clint_reset),
    .io_rtcTick(clint_io_rtcTick),
    .io_int_0_0(clint_io_int_0_0),
    .io_int_0_1(clint_io_int_0_1),
    .io_in_0_a_ready(clint_io_in_0_a_ready),
    .io_in_0_a_valid(clint_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(clint_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(clint_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(clint_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(clint_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(clint_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(clint_io_in_0_a_bits_data),
    .io_in_0_d_ready(clint_io_in_0_d_ready),
    .io_in_0_d_valid(clint_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(clint_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(clint_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(clint_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(clint_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(clint_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(clint_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(clint_io_in_0_d_bits_error)
  );
  TLDebugModule_debug debug_1 (
    .clock(debug_1_clock),
    .reset(debug_1_reset),
    .io_debugInterrupts_0_0(debug_1_io_debugInterrupts_0_0),
    .io_in_0_a_ready(debug_1_io_in_0_a_ready),
    .io_in_0_a_valid(debug_1_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(debug_1_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(debug_1_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(debug_1_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(debug_1_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(debug_1_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(debug_1_io_in_0_a_bits_data),
    .io_in_0_d_ready(debug_1_io_in_0_d_ready),
    .io_in_0_d_valid(debug_1_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(debug_1_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(debug_1_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(debug_1_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(debug_1_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(debug_1_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(debug_1_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(debug_1_io_in_0_d_bits_error),
    .io_ctrl_debugUnavail_0(debug_1_io_ctrl_debugUnavail_0),
    .io_ctrl_ndreset(debug_1_io_ctrl_ndreset),
    .io_dmi_dmi_req_ready(debug_1_io_dmi_dmi_req_ready),
    .io_dmi_dmi_req_valid(debug_1_io_dmi_dmi_req_valid),
    .io_dmi_dmi_req_bits_addr(debug_1_io_dmi_dmi_req_bits_addr),
    .io_dmi_dmi_req_bits_data(debug_1_io_dmi_dmi_req_bits_data),
    .io_dmi_dmi_req_bits_op(debug_1_io_dmi_dmi_req_bits_op),
    .io_dmi_dmi_resp_ready(debug_1_io_dmi_dmi_resp_ready),
    .io_dmi_dmi_resp_valid(debug_1_io_dmi_dmi_resp_valid),
    .io_dmi_dmi_resp_bits_data(debug_1_io_dmi_dmi_resp_bits_data),
    .io_dmi_dmi_resp_bits_resp(debug_1_io_dmi_dmi_resp_bits_resp),
    .io_dmi_dmiClock(debug_1_io_dmi_dmiClock),
    .io_dmi_dmiReset(debug_1_io_dmi_dmiReset)
  );
  SyncRocketTile_tile tile (
    .clock(tile_clock),
    .reset(tile_reset),
    .io_master_0_a_ready(tile_io_master_0_a_ready),
    .io_master_0_a_valid(tile_io_master_0_a_valid),
    .io_master_0_a_bits_opcode(tile_io_master_0_a_bits_opcode),
    .io_master_0_a_bits_param(tile_io_master_0_a_bits_param),
    .io_master_0_a_bits_size(tile_io_master_0_a_bits_size),
    .io_master_0_a_bits_source(tile_io_master_0_a_bits_source),
    .io_master_0_a_bits_address(tile_io_master_0_a_bits_address),
    .io_master_0_a_bits_mask(tile_io_master_0_a_bits_mask),
    .io_master_0_a_bits_data(tile_io_master_0_a_bits_data),
    .io_master_0_d_ready(tile_io_master_0_d_ready),
    .io_master_0_d_valid(tile_io_master_0_d_valid),
    .io_master_0_d_bits_opcode(tile_io_master_0_d_bits_opcode),
    .io_master_0_d_bits_size(tile_io_master_0_d_bits_size),
    .io_master_0_d_bits_source(tile_io_master_0_d_bits_source),
    .io_master_0_d_bits_data(tile_io_master_0_d_bits_data),
    .io_master_0_d_bits_error(tile_io_master_0_d_bits_error),
    .io_slave_0_a_ready(tile_io_slave_0_a_ready),
    .io_slave_0_a_valid(tile_io_slave_0_a_valid),
    .io_slave_0_a_bits_opcode(tile_io_slave_0_a_bits_opcode),
    .io_slave_0_a_bits_param(tile_io_slave_0_a_bits_param),
    .io_slave_0_a_bits_size(tile_io_slave_0_a_bits_size),
    .io_slave_0_a_bits_source(tile_io_slave_0_a_bits_source),
    .io_slave_0_a_bits_address(tile_io_slave_0_a_bits_address),
    .io_slave_0_a_bits_mask(tile_io_slave_0_a_bits_mask),
    .io_slave_0_a_bits_data(tile_io_slave_0_a_bits_data),
    .io_slave_0_d_ready(tile_io_slave_0_d_ready),
    .io_slave_0_d_valid(tile_io_slave_0_d_valid),
    .io_slave_0_d_bits_opcode(tile_io_slave_0_d_bits_opcode),
    .io_slave_0_d_bits_param(tile_io_slave_0_d_bits_param),
    .io_slave_0_d_bits_size(tile_io_slave_0_d_bits_size),
    .io_slave_0_d_bits_source(tile_io_slave_0_d_bits_source),
    .io_slave_0_d_bits_sink(tile_io_slave_0_d_bits_sink),
    .io_slave_0_d_bits_data(tile_io_slave_0_d_bits_data),
    .io_slave_0_d_bits_error(tile_io_slave_0_d_bits_error),
    .io_asyncInterrupts_0_0(tile_io_asyncInterrupts_0_0),
    .io_periphInterrupts_0_0(tile_io_periphInterrupts_0_0),
    .io_periphInterrupts_0_1(tile_io_periphInterrupts_0_1),
    .io_periphInterrupts_0_2(tile_io_periphInterrupts_0_2),
    .io_hartid(tile_io_hartid),
    .io_resetVector(tile_io_resetVector)
  );
  TLBuffer_4 TLBuffer_4 (
    .clock(TLBuffer_4_clock),
    .reset(TLBuffer_4_reset),
    .io_in_0_a_ready(TLBuffer_4_io_in_0_a_ready),
    .io_in_0_a_valid(TLBuffer_4_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLBuffer_4_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLBuffer_4_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLBuffer_4_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLBuffer_4_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLBuffer_4_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLBuffer_4_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLBuffer_4_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLBuffer_4_io_in_0_d_ready),
    .io_in_0_d_valid(TLBuffer_4_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLBuffer_4_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLBuffer_4_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLBuffer_4_io_in_0_d_bits_source),
    .io_in_0_d_bits_data(TLBuffer_4_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLBuffer_4_io_in_0_d_bits_error),
    .io_out_0_a_ready(TLBuffer_4_io_out_0_a_ready),
    .io_out_0_a_valid(TLBuffer_4_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLBuffer_4_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLBuffer_4_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLBuffer_4_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLBuffer_4_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLBuffer_4_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLBuffer_4_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLBuffer_4_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLBuffer_4_io_out_0_d_ready),
    .io_out_0_d_valid(TLBuffer_4_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLBuffer_4_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(TLBuffer_4_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLBuffer_4_io_out_0_d_bits_source),
    .io_out_0_d_bits_data(TLBuffer_4_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(TLBuffer_4_io_out_0_d_bits_error)
  );
  IntXbar_1 IntXbar_1 (
    .io_in_0_0(IntXbar_1_io_in_0_0),
    .io_out_0_0(IntXbar_1_io_out_0_0)
  );
  IntXbar_2 IntXbar_2 (
    .io_in_1_0(IntXbar_2_io_in_1_0),
    .io_in_0_0(IntXbar_2_io_in_0_0),
    .io_in_0_1(IntXbar_2_io_in_0_1),
    .io_out_0_0(IntXbar_2_io_out_0_0),
    .io_out_0_1(IntXbar_2_io_out_0_1),
    .io_out_0_2(IntXbar_2_io_out_0_2)
  );
  IntXing IntXing (
    .clock(IntXing_clock),
    .io_in_0_0(IntXing_io_in_0_0),
    .io_in_0_1(IntXing_io_in_0_1),
    .io_out_0_0(IntXing_io_out_0_0),
    .io_out_0_1(IntXing_io_out_0_1)
  );
  TLToAXI4 TLToAXI4 (
    .clock(TLToAXI4_clock),
    .reset(TLToAXI4_reset),
    .io_in_0_a_ready(TLToAXI4_io_in_0_a_ready),
    .io_in_0_a_valid(TLToAXI4_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLToAXI4_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(TLToAXI4_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLToAXI4_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLToAXI4_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLToAXI4_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLToAXI4_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLToAXI4_io_in_0_d_ready),
    .io_in_0_d_valid(TLToAXI4_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLToAXI4_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(TLToAXI4_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(TLToAXI4_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLToAXI4_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(TLToAXI4_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(TLToAXI4_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(TLToAXI4_io_in_0_d_bits_error),
    .io_out_0_aw_ready(TLToAXI4_io_out_0_aw_ready),
    .io_out_0_aw_valid(TLToAXI4_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(TLToAXI4_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(TLToAXI4_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(TLToAXI4_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(TLToAXI4_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_burst(TLToAXI4_io_out_0_aw_bits_burst),
    .io_out_0_aw_bits_user(TLToAXI4_io_out_0_aw_bits_user),
    .io_out_0_w_ready(TLToAXI4_io_out_0_w_ready),
    .io_out_0_w_valid(TLToAXI4_io_out_0_w_valid),
    .io_out_0_w_bits_data(TLToAXI4_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(TLToAXI4_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(TLToAXI4_io_out_0_w_bits_last),
    .io_out_0_b_ready(TLToAXI4_io_out_0_b_ready),
    .io_out_0_b_valid(TLToAXI4_io_out_0_b_valid),
    .io_out_0_b_bits_id(TLToAXI4_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(TLToAXI4_io_out_0_b_bits_resp),
    .io_out_0_b_bits_user(TLToAXI4_io_out_0_b_bits_user),
    .io_out_0_ar_ready(TLToAXI4_io_out_0_ar_ready),
    .io_out_0_ar_valid(TLToAXI4_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(TLToAXI4_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(TLToAXI4_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(TLToAXI4_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(TLToAXI4_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_burst(TLToAXI4_io_out_0_ar_bits_burst),
    .io_out_0_ar_bits_user(TLToAXI4_io_out_0_ar_bits_user),
    .io_out_0_r_ready(TLToAXI4_io_out_0_r_ready),
    .io_out_0_r_valid(TLToAXI4_io_out_0_r_valid),
    .io_out_0_r_bits_id(TLToAXI4_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(TLToAXI4_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(TLToAXI4_io_out_0_r_bits_resp),
    .io_out_0_r_bits_user(TLToAXI4_io_out_0_r_bits_user),
    .io_out_0_r_bits_last(TLToAXI4_io_out_0_r_bits_last)
  );
  AXI4IdIndexer AXI4IdIndexer (
    .io_in_0_aw_ready(AXI4IdIndexer_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4IdIndexer_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4IdIndexer_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4IdIndexer_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4IdIndexer_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4IdIndexer_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4IdIndexer_io_in_0_aw_bits_burst),
    .io_in_0_aw_bits_user(AXI4IdIndexer_io_in_0_aw_bits_user),
    .io_in_0_w_ready(AXI4IdIndexer_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4IdIndexer_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4IdIndexer_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4IdIndexer_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4IdIndexer_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4IdIndexer_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4IdIndexer_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4IdIndexer_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4IdIndexer_io_in_0_b_bits_resp),
    .io_in_0_b_bits_user(AXI4IdIndexer_io_in_0_b_bits_user),
    .io_in_0_ar_ready(AXI4IdIndexer_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4IdIndexer_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4IdIndexer_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4IdIndexer_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4IdIndexer_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4IdIndexer_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4IdIndexer_io_in_0_ar_bits_burst),
    .io_in_0_ar_bits_user(AXI4IdIndexer_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4IdIndexer_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4IdIndexer_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4IdIndexer_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4IdIndexer_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4IdIndexer_io_in_0_r_bits_resp),
    .io_in_0_r_bits_user(AXI4IdIndexer_io_in_0_r_bits_user),
    .io_in_0_r_bits_last(AXI4IdIndexer_io_in_0_r_bits_last),
    .io_out_0_aw_ready(AXI4IdIndexer_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4IdIndexer_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4IdIndexer_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4IdIndexer_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4IdIndexer_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4IdIndexer_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_burst(AXI4IdIndexer_io_out_0_aw_bits_burst),
    .io_out_0_aw_bits_user(AXI4IdIndexer_io_out_0_aw_bits_user),
    .io_out_0_w_ready(AXI4IdIndexer_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4IdIndexer_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4IdIndexer_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4IdIndexer_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4IdIndexer_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4IdIndexer_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4IdIndexer_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4IdIndexer_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(AXI4IdIndexer_io_out_0_b_bits_resp),
    .io_out_0_b_bits_user(AXI4IdIndexer_io_out_0_b_bits_user),
    .io_out_0_ar_ready(AXI4IdIndexer_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4IdIndexer_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4IdIndexer_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4IdIndexer_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4IdIndexer_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4IdIndexer_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_burst(AXI4IdIndexer_io_out_0_ar_bits_burst),
    .io_out_0_ar_bits_user(AXI4IdIndexer_io_out_0_ar_bits_user),
    .io_out_0_r_ready(AXI4IdIndexer_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4IdIndexer_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4IdIndexer_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(AXI4IdIndexer_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(AXI4IdIndexer_io_out_0_r_bits_resp),
    .io_out_0_r_bits_user(AXI4IdIndexer_io_out_0_r_bits_user),
    .io_out_0_r_bits_last(AXI4IdIndexer_io_out_0_r_bits_last)
  );
  AXI4Deinterleaver AXI4Deinterleaver (
    .clock(AXI4Deinterleaver_clock),
    .reset(AXI4Deinterleaver_reset),
    .io_in_0_aw_ready(AXI4Deinterleaver_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4Deinterleaver_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4Deinterleaver_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4Deinterleaver_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4Deinterleaver_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4Deinterleaver_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4Deinterleaver_io_in_0_aw_bits_burst),
    .io_in_0_aw_bits_user(AXI4Deinterleaver_io_in_0_aw_bits_user),
    .io_in_0_w_ready(AXI4Deinterleaver_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4Deinterleaver_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4Deinterleaver_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4Deinterleaver_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4Deinterleaver_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4Deinterleaver_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4Deinterleaver_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4Deinterleaver_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4Deinterleaver_io_in_0_b_bits_resp),
    .io_in_0_b_bits_user(AXI4Deinterleaver_io_in_0_b_bits_user),
    .io_in_0_ar_ready(AXI4Deinterleaver_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4Deinterleaver_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4Deinterleaver_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4Deinterleaver_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4Deinterleaver_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4Deinterleaver_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4Deinterleaver_io_in_0_ar_bits_burst),
    .io_in_0_ar_bits_user(AXI4Deinterleaver_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4Deinterleaver_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4Deinterleaver_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4Deinterleaver_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4Deinterleaver_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4Deinterleaver_io_in_0_r_bits_resp),
    .io_in_0_r_bits_user(AXI4Deinterleaver_io_in_0_r_bits_user),
    .io_in_0_r_bits_last(AXI4Deinterleaver_io_in_0_r_bits_last),
    .io_out_0_aw_ready(AXI4Deinterleaver_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4Deinterleaver_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4Deinterleaver_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4Deinterleaver_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4Deinterleaver_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4Deinterleaver_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_burst(AXI4Deinterleaver_io_out_0_aw_bits_burst),
    .io_out_0_aw_bits_user(AXI4Deinterleaver_io_out_0_aw_bits_user),
    .io_out_0_w_ready(AXI4Deinterleaver_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4Deinterleaver_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4Deinterleaver_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4Deinterleaver_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4Deinterleaver_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4Deinterleaver_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4Deinterleaver_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4Deinterleaver_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(AXI4Deinterleaver_io_out_0_b_bits_resp),
    .io_out_0_b_bits_user(AXI4Deinterleaver_io_out_0_b_bits_user),
    .io_out_0_ar_ready(AXI4Deinterleaver_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4Deinterleaver_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4Deinterleaver_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4Deinterleaver_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4Deinterleaver_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4Deinterleaver_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_burst(AXI4Deinterleaver_io_out_0_ar_bits_burst),
    .io_out_0_ar_bits_user(AXI4Deinterleaver_io_out_0_ar_bits_user),
    .io_out_0_r_ready(AXI4Deinterleaver_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4Deinterleaver_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4Deinterleaver_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(AXI4Deinterleaver_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(AXI4Deinterleaver_io_out_0_r_bits_resp),
    .io_out_0_r_bits_user(AXI4Deinterleaver_io_out_0_r_bits_user),
    .io_out_0_r_bits_last(AXI4Deinterleaver_io_out_0_r_bits_last)
  );
  AXI4UserYanker AXI4UserYanker (
    .clock(AXI4UserYanker_clock),
    .reset(AXI4UserYanker_reset),
    .io_in_0_aw_ready(AXI4UserYanker_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4UserYanker_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4UserYanker_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4UserYanker_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4UserYanker_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4UserYanker_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4UserYanker_io_in_0_aw_bits_burst),
    .io_in_0_aw_bits_user(AXI4UserYanker_io_in_0_aw_bits_user),
    .io_in_0_w_ready(AXI4UserYanker_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4UserYanker_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4UserYanker_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4UserYanker_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4UserYanker_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4UserYanker_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4UserYanker_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4UserYanker_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4UserYanker_io_in_0_b_bits_resp),
    .io_in_0_b_bits_user(AXI4UserYanker_io_in_0_b_bits_user),
    .io_in_0_ar_ready(AXI4UserYanker_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4UserYanker_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4UserYanker_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4UserYanker_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4UserYanker_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4UserYanker_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4UserYanker_io_in_0_ar_bits_burst),
    .io_in_0_ar_bits_user(AXI4UserYanker_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4UserYanker_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4UserYanker_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4UserYanker_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4UserYanker_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4UserYanker_io_in_0_r_bits_resp),
    .io_in_0_r_bits_user(AXI4UserYanker_io_in_0_r_bits_user),
    .io_in_0_r_bits_last(AXI4UserYanker_io_in_0_r_bits_last),
    .io_out_0_aw_ready(AXI4UserYanker_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4UserYanker_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4UserYanker_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4UserYanker_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4UserYanker_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4UserYanker_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_burst(AXI4UserYanker_io_out_0_aw_bits_burst),
    .io_out_0_w_ready(AXI4UserYanker_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4UserYanker_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4UserYanker_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4UserYanker_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4UserYanker_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4UserYanker_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4UserYanker_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4UserYanker_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(AXI4UserYanker_io_out_0_b_bits_resp),
    .io_out_0_ar_ready(AXI4UserYanker_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4UserYanker_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4UserYanker_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4UserYanker_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4UserYanker_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4UserYanker_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_burst(AXI4UserYanker_io_out_0_ar_bits_burst),
    .io_out_0_r_ready(AXI4UserYanker_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4UserYanker_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4UserYanker_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(AXI4UserYanker_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(AXI4UserYanker_io_out_0_r_bits_resp),
    .io_out_0_r_bits_last(AXI4UserYanker_io_out_0_r_bits_last)
  );
  AXI4Buffer AXI4Buffer (
    .clock(AXI4Buffer_clock),
    .reset(AXI4Buffer_reset),
    .io_in_0_aw_ready(AXI4Buffer_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4Buffer_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4Buffer_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4Buffer_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4Buffer_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4Buffer_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4Buffer_io_in_0_aw_bits_burst),
    .io_in_0_w_ready(AXI4Buffer_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4Buffer_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4Buffer_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4Buffer_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4Buffer_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4Buffer_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4Buffer_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4Buffer_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4Buffer_io_in_0_b_bits_resp),
    .io_in_0_ar_ready(AXI4Buffer_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4Buffer_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4Buffer_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4Buffer_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4Buffer_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4Buffer_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4Buffer_io_in_0_ar_bits_burst),
    .io_in_0_r_ready(AXI4Buffer_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4Buffer_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4Buffer_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4Buffer_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4Buffer_io_in_0_r_bits_resp),
    .io_in_0_r_bits_last(AXI4Buffer_io_in_0_r_bits_last),
    .io_out_0_aw_ready(AXI4Buffer_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4Buffer_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4Buffer_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4Buffer_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4Buffer_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4Buffer_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_burst(AXI4Buffer_io_out_0_aw_bits_burst),
    .io_out_0_w_ready(AXI4Buffer_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4Buffer_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4Buffer_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4Buffer_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4Buffer_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4Buffer_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4Buffer_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4Buffer_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(AXI4Buffer_io_out_0_b_bits_resp),
    .io_out_0_ar_ready(AXI4Buffer_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4Buffer_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4Buffer_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4Buffer_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4Buffer_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4Buffer_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_burst(AXI4Buffer_io_out_0_ar_bits_burst),
    .io_out_0_r_ready(AXI4Buffer_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4Buffer_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4Buffer_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(AXI4Buffer_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(AXI4Buffer_io_out_0_r_bits_resp),
    .io_out_0_r_bits_last(AXI4Buffer_io_out_0_r_bits_last)
  );
  TLBuffer_5 TLBuffer_5 (
    .clock(TLBuffer_5_clock),
    .reset(TLBuffer_5_reset),
    .io_in_0_a_ready(TLBuffer_5_io_in_0_a_ready),
    .io_in_0_a_valid(TLBuffer_5_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLBuffer_5_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLBuffer_5_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLBuffer_5_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLBuffer_5_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLBuffer_5_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLBuffer_5_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLBuffer_5_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLBuffer_5_io_in_0_d_ready),
    .io_in_0_d_valid(TLBuffer_5_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLBuffer_5_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLBuffer_5_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLBuffer_5_io_in_0_d_bits_source),
    .io_out_0_a_ready(TLBuffer_5_io_out_0_a_ready),
    .io_out_0_a_valid(TLBuffer_5_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLBuffer_5_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLBuffer_5_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLBuffer_5_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLBuffer_5_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLBuffer_5_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLBuffer_5_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLBuffer_5_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLBuffer_5_io_out_0_d_ready),
    .io_out_0_d_valid(TLBuffer_5_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLBuffer_5_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(TLBuffer_5_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLBuffer_5_io_out_0_d_bits_source)
  );
  AXI4IdIndexer_1 AXI4IdIndexer_1 (
    .io_in_0_aw_valid(AXI4IdIndexer_1_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4IdIndexer_1_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4IdIndexer_1_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4IdIndexer_1_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4IdIndexer_1_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4IdIndexer_1_io_in_0_aw_bits_burst),
    .io_in_0_w_valid(AXI4IdIndexer_1_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4IdIndexer_1_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4IdIndexer_1_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4IdIndexer_1_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4IdIndexer_1_io_in_0_b_ready),
    .io_in_0_ar_valid(AXI4IdIndexer_1_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4IdIndexer_1_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4IdIndexer_1_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4IdIndexer_1_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4IdIndexer_1_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4IdIndexer_1_io_in_0_ar_bits_burst),
    .io_in_0_r_ready(AXI4IdIndexer_1_io_in_0_r_ready),
    .io_out_0_aw_valid(AXI4IdIndexer_1_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4IdIndexer_1_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4IdIndexer_1_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4IdIndexer_1_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4IdIndexer_1_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_burst(AXI4IdIndexer_1_io_out_0_aw_bits_burst),
    .io_out_0_aw_bits_user(AXI4IdIndexer_1_io_out_0_aw_bits_user),
    .io_out_0_w_valid(AXI4IdIndexer_1_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4IdIndexer_1_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4IdIndexer_1_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4IdIndexer_1_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4IdIndexer_1_io_out_0_b_ready),
    .io_out_0_ar_valid(AXI4IdIndexer_1_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4IdIndexer_1_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4IdIndexer_1_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4IdIndexer_1_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4IdIndexer_1_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_burst(AXI4IdIndexer_1_io_out_0_ar_bits_burst),
    .io_out_0_ar_bits_user(AXI4IdIndexer_1_io_out_0_ar_bits_user),
    .io_out_0_r_ready(AXI4IdIndexer_1_io_out_0_r_ready)
  );
  AXI4Fragmenter AXI4Fragmenter (
    .clock(AXI4Fragmenter_clock),
    .reset(AXI4Fragmenter_reset),
    .io_in_0_aw_valid(AXI4Fragmenter_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4Fragmenter_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4Fragmenter_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4Fragmenter_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4Fragmenter_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4Fragmenter_io_in_0_aw_bits_burst),
    .io_in_0_aw_bits_user(AXI4Fragmenter_io_in_0_aw_bits_user),
    .io_in_0_w_valid(AXI4Fragmenter_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4Fragmenter_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4Fragmenter_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4Fragmenter_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4Fragmenter_io_in_0_b_ready),
    .io_in_0_ar_valid(AXI4Fragmenter_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4Fragmenter_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4Fragmenter_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4Fragmenter_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4Fragmenter_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4Fragmenter_io_in_0_ar_bits_burst),
    .io_in_0_ar_bits_user(AXI4Fragmenter_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4Fragmenter_io_in_0_r_ready),
    .io_out_0_aw_ready(AXI4Fragmenter_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4Fragmenter_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4Fragmenter_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4Fragmenter_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4Fragmenter_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4Fragmenter_io_out_0_aw_bits_size),
    .io_out_0_aw_bits_user(AXI4Fragmenter_io_out_0_aw_bits_user),
    .io_out_0_w_ready(AXI4Fragmenter_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4Fragmenter_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4Fragmenter_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4Fragmenter_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4Fragmenter_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4Fragmenter_io_out_0_b_ready),
    .io_out_0_b_bits_user(AXI4Fragmenter_io_out_0_b_bits_user),
    .io_out_0_ar_ready(AXI4Fragmenter_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4Fragmenter_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4Fragmenter_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4Fragmenter_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4Fragmenter_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4Fragmenter_io_out_0_ar_bits_size),
    .io_out_0_ar_bits_user(AXI4Fragmenter_io_out_0_ar_bits_user),
    .io_out_0_r_ready(AXI4Fragmenter_io_out_0_r_ready)
  );
  AXI4UserYanker_1 AXI4UserYanker_1 (
    .clock(AXI4UserYanker_1_clock),
    .reset(AXI4UserYanker_1_reset),
    .io_in_0_aw_ready(AXI4UserYanker_1_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4UserYanker_1_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4UserYanker_1_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4UserYanker_1_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4UserYanker_1_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4UserYanker_1_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_user(AXI4UserYanker_1_io_in_0_aw_bits_user),
    .io_in_0_w_ready(AXI4UserYanker_1_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4UserYanker_1_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4UserYanker_1_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4UserYanker_1_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4UserYanker_1_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4UserYanker_1_io_in_0_b_ready),
    .io_in_0_b_bits_user(AXI4UserYanker_1_io_in_0_b_bits_user),
    .io_in_0_ar_ready(AXI4UserYanker_1_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4UserYanker_1_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4UserYanker_1_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4UserYanker_1_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4UserYanker_1_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4UserYanker_1_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_user(AXI4UserYanker_1_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4UserYanker_1_io_in_0_r_ready),
    .io_out_0_aw_ready(AXI4UserYanker_1_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4UserYanker_1_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4UserYanker_1_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4UserYanker_1_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_len(AXI4UserYanker_1_io_out_0_aw_bits_len),
    .io_out_0_aw_bits_size(AXI4UserYanker_1_io_out_0_aw_bits_size),
    .io_out_0_w_ready(AXI4UserYanker_1_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4UserYanker_1_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4UserYanker_1_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4UserYanker_1_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4UserYanker_1_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4UserYanker_1_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4UserYanker_1_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4UserYanker_1_io_out_0_b_bits_id),
    .io_out_0_ar_ready(AXI4UserYanker_1_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4UserYanker_1_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4UserYanker_1_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4UserYanker_1_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_len(AXI4UserYanker_1_io_out_0_ar_bits_len),
    .io_out_0_ar_bits_size(AXI4UserYanker_1_io_out_0_ar_bits_size),
    .io_out_0_r_ready(AXI4UserYanker_1_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4UserYanker_1_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4UserYanker_1_io_out_0_r_bits_id),
    .io_out_0_r_bits_last(AXI4UserYanker_1_io_out_0_r_bits_last)
  );
  AXI4ToTL AXI4ToTL (
    .clock(AXI4ToTL_clock),
    .reset(AXI4ToTL_reset),
    .io_in_0_aw_ready(AXI4ToTL_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4ToTL_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4ToTL_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4ToTL_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4ToTL_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4ToTL_io_in_0_aw_bits_size),
    .io_in_0_w_ready(AXI4ToTL_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4ToTL_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4ToTL_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4ToTL_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4ToTL_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4ToTL_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4ToTL_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4ToTL_io_in_0_b_bits_id),
    .io_in_0_ar_ready(AXI4ToTL_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4ToTL_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4ToTL_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4ToTL_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4ToTL_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4ToTL_io_in_0_ar_bits_size),
    .io_in_0_r_ready(AXI4ToTL_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4ToTL_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4ToTL_io_in_0_r_bits_id),
    .io_in_0_r_bits_last(AXI4ToTL_io_in_0_r_bits_last),
    .io_out_0_a_ready(AXI4ToTL_io_out_0_a_ready),
    .io_out_0_a_valid(AXI4ToTL_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(AXI4ToTL_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(AXI4ToTL_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(AXI4ToTL_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(AXI4ToTL_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(AXI4ToTL_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(AXI4ToTL_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(AXI4ToTL_io_out_0_a_bits_data),
    .io_out_0_d_ready(AXI4ToTL_io_out_0_d_ready),
    .io_out_0_d_valid(AXI4ToTL_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(AXI4ToTL_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(AXI4ToTL_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(AXI4ToTL_io_out_0_d_bits_source)
  );
  TLWidthWidget_2 TLWidthWidget_2 (
    .clock(TLWidthWidget_2_clock),
    .reset(TLWidthWidget_2_reset),
    .io_in_0_a_ready(TLWidthWidget_2_io_in_0_a_ready),
    .io_in_0_a_valid(TLWidthWidget_2_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(TLWidthWidget_2_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_param(TLWidthWidget_2_io_in_0_a_bits_param),
    .io_in_0_a_bits_size(TLWidthWidget_2_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(TLWidthWidget_2_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(TLWidthWidget_2_io_in_0_a_bits_address),
    .io_in_0_a_bits_mask(TLWidthWidget_2_io_in_0_a_bits_mask),
    .io_in_0_a_bits_data(TLWidthWidget_2_io_in_0_a_bits_data),
    .io_in_0_d_ready(TLWidthWidget_2_io_in_0_d_ready),
    .io_in_0_d_valid(TLWidthWidget_2_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(TLWidthWidget_2_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_size(TLWidthWidget_2_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(TLWidthWidget_2_io_in_0_d_bits_source),
    .io_out_0_a_ready(TLWidthWidget_2_io_out_0_a_ready),
    .io_out_0_a_valid(TLWidthWidget_2_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(TLWidthWidget_2_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_param(TLWidthWidget_2_io_out_0_a_bits_param),
    .io_out_0_a_bits_size(TLWidthWidget_2_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(TLWidthWidget_2_io_out_0_a_bits_source),
    .io_out_0_a_bits_address(TLWidthWidget_2_io_out_0_a_bits_address),
    .io_out_0_a_bits_mask(TLWidthWidget_2_io_out_0_a_bits_mask),
    .io_out_0_a_bits_data(TLWidthWidget_2_io_out_0_a_bits_data),
    .io_out_0_d_ready(TLWidthWidget_2_io_out_0_d_ready),
    .io_out_0_d_valid(TLWidthWidget_2_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(TLWidthWidget_2_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_size(TLWidthWidget_2_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(TLWidthWidget_2_io_out_0_d_bits_source)
  );
  TLROM_bootrom bootrom (
    .io_in_0_a_ready(bootrom_io_in_0_a_ready),
    .io_in_0_a_valid(bootrom_io_in_0_a_valid),
    .io_in_0_a_bits_size(bootrom_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(bootrom_io_in_0_a_bits_source),
    .io_in_0_a_bits_address(bootrom_io_in_0_a_bits_address),
    .io_in_0_d_ready(bootrom_io_in_0_d_ready),
    .io_in_0_d_valid(bootrom_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(bootrom_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(bootrom_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(bootrom_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(bootrom_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(bootrom_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(bootrom_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(bootrom_io_in_0_d_bits_error)
  );
  TLError_error error (
    .clock(error_clock),
    .reset(error_reset),
    .io_in_0_a_ready(error_io_in_0_a_ready),
    .io_in_0_a_valid(error_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(error_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(error_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(error_io_in_0_a_bits_source),
    .io_in_0_c_valid(error_io_in_0_c_valid),
    .io_in_0_c_bits_param(error_io_in_0_c_bits_param),
    .io_in_0_c_bits_size(error_io_in_0_c_bits_size),
    .io_in_0_c_bits_source(error_io_in_0_c_bits_source),
    .io_in_0_d_ready(error_io_in_0_d_ready),
    .io_in_0_d_valid(error_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(error_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(error_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(error_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(error_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(error_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(error_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(error_io_in_0_d_bits_error)
  );
  TLBuffer_error error_TLBuffer (
    .clock(error_TLBuffer_clock),
    .reset(error_TLBuffer_reset),
    .io_in_0_a_ready(error_TLBuffer_io_in_0_a_ready),
    .io_in_0_a_valid(error_TLBuffer_io_in_0_a_valid),
    .io_in_0_a_bits_opcode(error_TLBuffer_io_in_0_a_bits_opcode),
    .io_in_0_a_bits_size(error_TLBuffer_io_in_0_a_bits_size),
    .io_in_0_a_bits_source(error_TLBuffer_io_in_0_a_bits_source),
    .io_in_0_d_ready(error_TLBuffer_io_in_0_d_ready),
    .io_in_0_d_valid(error_TLBuffer_io_in_0_d_valid),
    .io_in_0_d_bits_opcode(error_TLBuffer_io_in_0_d_bits_opcode),
    .io_in_0_d_bits_param(error_TLBuffer_io_in_0_d_bits_param),
    .io_in_0_d_bits_size(error_TLBuffer_io_in_0_d_bits_size),
    .io_in_0_d_bits_source(error_TLBuffer_io_in_0_d_bits_source),
    .io_in_0_d_bits_sink(error_TLBuffer_io_in_0_d_bits_sink),
    .io_in_0_d_bits_data(error_TLBuffer_io_in_0_d_bits_data),
    .io_in_0_d_bits_error(error_TLBuffer_io_in_0_d_bits_error),
    .io_out_0_a_ready(error_TLBuffer_io_out_0_a_ready),
    .io_out_0_a_valid(error_TLBuffer_io_out_0_a_valid),
    .io_out_0_a_bits_opcode(error_TLBuffer_io_out_0_a_bits_opcode),
    .io_out_0_a_bits_size(error_TLBuffer_io_out_0_a_bits_size),
    .io_out_0_a_bits_source(error_TLBuffer_io_out_0_a_bits_source),
    .io_out_0_c_valid(error_TLBuffer_io_out_0_c_valid),
    .io_out_0_c_bits_param(error_TLBuffer_io_out_0_c_bits_param),
    .io_out_0_c_bits_size(error_TLBuffer_io_out_0_c_bits_size),
    .io_out_0_c_bits_source(error_TLBuffer_io_out_0_c_bits_source),
    .io_out_0_d_ready(error_TLBuffer_io_out_0_d_ready),
    .io_out_0_d_valid(error_TLBuffer_io_out_0_d_valid),
    .io_out_0_d_bits_opcode(error_TLBuffer_io_out_0_d_bits_opcode),
    .io_out_0_d_bits_param(error_TLBuffer_io_out_0_d_bits_param),
    .io_out_0_d_bits_size(error_TLBuffer_io_out_0_d_bits_size),
    .io_out_0_d_bits_source(error_TLBuffer_io_out_0_d_bits_source),
    .io_out_0_d_bits_sink(error_TLBuffer_io_out_0_d_bits_sink),
    .io_out_0_d_bits_data(error_TLBuffer_io_out_0_d_bits_data),
    .io_out_0_d_bits_error(error_TLBuffer_io_out_0_d_bits_error)
  );
  assign debug_clockeddmi_dmi_req_ready = debug_1_io_dmi_dmi_req_ready;
  assign debug_clockeddmi_dmi_resp_valid = debug_1_io_dmi_dmi_resp_valid;
  assign debug_clockeddmi_dmi_resp_bits_data = debug_1_io_dmi_dmi_resp_bits_data;
  assign debug_clockeddmi_dmi_resp_bits_resp = debug_1_io_dmi_dmi_resp_bits_resp;
  assign debug_ndreset = debug_1_io_ctrl_ndreset;
  assign mmio_axi4_0_aw_valid = AXI4Buffer_io_out_0_aw_valid;
  assign mmio_axi4_0_aw_bits_id = AXI4Buffer_io_out_0_aw_bits_id;
  assign mmio_axi4_0_aw_bits_addr = AXI4Buffer_io_out_0_aw_bits_addr;
  assign mmio_axi4_0_aw_bits_len = AXI4Buffer_io_out_0_aw_bits_len;
  assign mmio_axi4_0_aw_bits_size = AXI4Buffer_io_out_0_aw_bits_size;
  assign mmio_axi4_0_aw_bits_burst = AXI4Buffer_io_out_0_aw_bits_burst;
  assign mmio_axi4_0_w_valid = AXI4Buffer_io_out_0_w_valid;
  assign mmio_axi4_0_w_bits_data = AXI4Buffer_io_out_0_w_bits_data;
  assign mmio_axi4_0_w_bits_strb = AXI4Buffer_io_out_0_w_bits_strb;
  assign mmio_axi4_0_w_bits_last = AXI4Buffer_io_out_0_w_bits_last;
  assign mmio_axi4_0_b_ready = AXI4Buffer_io_out_0_b_ready;
  assign mmio_axi4_0_ar_valid = AXI4Buffer_io_out_0_ar_valid;
  assign mmio_axi4_0_ar_bits_id = AXI4Buffer_io_out_0_ar_bits_id;
  assign mmio_axi4_0_ar_bits_addr = AXI4Buffer_io_out_0_ar_bits_addr;
  assign mmio_axi4_0_ar_bits_len = AXI4Buffer_io_out_0_ar_bits_len;
  assign mmio_axi4_0_ar_bits_size = AXI4Buffer_io_out_0_ar_bits_size;
  assign mmio_axi4_0_ar_bits_burst = AXI4Buffer_io_out_0_ar_bits_burst;
  assign mmio_axi4_0_r_ready = AXI4Buffer_io_out_0_r_ready;
  assign IntXbar_io_in_0_0 = IntXing_io_out_0_0;
  assign IntXbar_io_in_0_1 = IntXing_io_out_0_1;
  assign TLXbar_clock = clock;
  assign TLXbar_reset = reset;
  assign TLXbar_io_in_1_a_valid = TLSplitter_io_out_1_a_valid;
  assign TLXbar_io_in_1_a_bits_opcode = TLSplitter_io_out_1_a_bits_opcode;
  assign TLXbar_io_in_1_a_bits_param = TLSplitter_io_out_1_a_bits_param;
  assign TLXbar_io_in_1_a_bits_size = TLSplitter_io_out_1_a_bits_size;
  assign TLXbar_io_in_1_a_bits_source = TLSplitter_io_out_1_a_bits_source;
  assign TLXbar_io_in_1_a_bits_address = TLSplitter_io_out_1_a_bits_address;
  assign TLXbar_io_in_1_a_bits_mask = TLSplitter_io_out_1_a_bits_mask;
  assign TLXbar_io_in_1_a_bits_data = TLSplitter_io_out_1_a_bits_data;
  assign TLXbar_io_in_1_d_ready = TLSplitter_io_out_1_d_ready;
  assign TLXbar_io_in_0_a_valid = TLSplitter_io_out_0_a_valid;
  assign TLXbar_io_in_0_a_bits_opcode = TLSplitter_io_out_0_a_bits_opcode;
  assign TLXbar_io_in_0_a_bits_param = TLSplitter_io_out_0_a_bits_param;
  assign TLXbar_io_in_0_a_bits_size = TLSplitter_io_out_0_a_bits_size;
  assign TLXbar_io_in_0_a_bits_source = TLSplitter_io_out_0_a_bits_source;
  assign TLXbar_io_in_0_a_bits_address = TLSplitter_io_out_0_a_bits_address;
  assign TLXbar_io_in_0_a_bits_mask = TLSplitter_io_out_0_a_bits_mask;
  assign TLXbar_io_in_0_a_bits_data = TLSplitter_io_out_0_a_bits_data;
  assign TLXbar_io_in_0_d_ready = TLSplitter_io_out_0_d_ready;
  assign TLXbar_io_out_2_a_ready = TLBuffer_1_io_in_2_a_ready;
  assign TLXbar_io_out_2_d_valid = TLBuffer_1_io_in_2_d_valid;
  assign TLXbar_io_out_2_d_bits_opcode = TLBuffer_1_io_in_2_d_bits_opcode;
  assign TLXbar_io_out_2_d_bits_param = TLBuffer_1_io_in_2_d_bits_param;
  assign TLXbar_io_out_2_d_bits_size = TLBuffer_1_io_in_2_d_bits_size;
  assign TLXbar_io_out_2_d_bits_source = TLBuffer_1_io_in_2_d_bits_source;
  assign TLXbar_io_out_2_d_bits_sink = TLBuffer_1_io_in_2_d_bits_sink;
  assign TLXbar_io_out_2_d_bits_data = TLBuffer_1_io_in_2_d_bits_data;
  assign TLXbar_io_out_2_d_bits_error = TLBuffer_1_io_in_2_d_bits_error;
  assign TLXbar_io_out_1_a_ready = TLBuffer_1_io_in_1_a_ready;
  assign TLXbar_io_out_1_d_valid = TLBuffer_1_io_in_1_d_valid;
  assign TLXbar_io_out_1_d_bits_opcode = TLBuffer_1_io_in_1_d_bits_opcode;
  assign TLXbar_io_out_1_d_bits_param = TLBuffer_1_io_in_1_d_bits_param;
  assign TLXbar_io_out_1_d_bits_size = TLBuffer_1_io_in_1_d_bits_size;
  assign TLXbar_io_out_1_d_bits_source = TLBuffer_1_io_in_1_d_bits_source;
  assign TLXbar_io_out_1_d_bits_sink = TLBuffer_1_io_in_1_d_bits_sink;
  assign TLXbar_io_out_1_d_bits_data = TLBuffer_1_io_in_1_d_bits_data;
  assign TLXbar_io_out_1_d_bits_error = TLBuffer_1_io_in_1_d_bits_error;
  assign TLXbar_io_out_0_a_ready = TLBuffer_1_io_in_0_a_ready;
  assign TLXbar_io_out_0_d_valid = TLBuffer_1_io_in_0_d_valid;
  assign TLXbar_io_out_0_d_bits_opcode = TLBuffer_1_io_in_0_d_bits_opcode;
  assign TLXbar_io_out_0_d_bits_param = TLBuffer_1_io_in_0_d_bits_param;
  assign TLXbar_io_out_0_d_bits_size = TLBuffer_1_io_in_0_d_bits_size;
  assign TLXbar_io_out_0_d_bits_source = TLBuffer_1_io_in_0_d_bits_source;
  assign TLXbar_io_out_0_d_bits_sink = TLBuffer_1_io_in_0_d_bits_sink;
  assign TLXbar_io_out_0_d_bits_data = TLBuffer_1_io_in_0_d_bits_data;
  assign TLXbar_io_out_0_d_bits_error = TLBuffer_1_io_in_0_d_bits_error;
  assign TLBuffer_1_clock = clock;
  assign TLBuffer_1_reset = reset;
  assign TLBuffer_1_io_in_2_a_valid = TLXbar_io_out_2_a_valid;
  assign TLBuffer_1_io_in_2_a_bits_opcode = TLXbar_io_out_2_a_bits_opcode;
  assign TLBuffer_1_io_in_2_a_bits_size = TLXbar_io_out_2_a_bits_size;
  assign TLBuffer_1_io_in_2_a_bits_source = TLXbar_io_out_2_a_bits_source;
  assign TLBuffer_1_io_in_2_d_ready = TLXbar_io_out_2_d_ready;
  assign TLBuffer_1_io_in_1_a_valid = TLXbar_io_out_1_a_valid;
  assign TLBuffer_1_io_in_1_a_bits_opcode = TLXbar_io_out_1_a_bits_opcode;
  assign TLBuffer_1_io_in_1_a_bits_size = TLXbar_io_out_1_a_bits_size;
  assign TLBuffer_1_io_in_1_a_bits_source = TLXbar_io_out_1_a_bits_source;
  assign TLBuffer_1_io_in_1_a_bits_address = TLXbar_io_out_1_a_bits_address;
  assign TLBuffer_1_io_in_1_a_bits_mask = TLXbar_io_out_1_a_bits_mask;
  assign TLBuffer_1_io_in_1_a_bits_data = TLXbar_io_out_1_a_bits_data;
  assign TLBuffer_1_io_in_1_d_ready = TLXbar_io_out_1_d_ready;
  assign TLBuffer_1_io_in_0_a_valid = TLXbar_io_out_0_a_valid;
  assign TLBuffer_1_io_in_0_a_bits_opcode = TLXbar_io_out_0_a_bits_opcode;
  assign TLBuffer_1_io_in_0_a_bits_param = TLXbar_io_out_0_a_bits_param;
  assign TLBuffer_1_io_in_0_a_bits_size = TLXbar_io_out_0_a_bits_size;
  assign TLBuffer_1_io_in_0_a_bits_source = TLXbar_io_out_0_a_bits_source;
  assign TLBuffer_1_io_in_0_a_bits_address = TLXbar_io_out_0_a_bits_address;
  assign TLBuffer_1_io_in_0_a_bits_mask = TLXbar_io_out_0_a_bits_mask;
  assign TLBuffer_1_io_in_0_a_bits_data = TLXbar_io_out_0_a_bits_data;
  assign TLBuffer_1_io_in_0_d_ready = TLXbar_io_out_0_d_ready;
  assign TLBuffer_1_io_out_2_a_ready = error_TLBuffer_io_in_0_a_ready;
  assign TLBuffer_1_io_out_2_d_valid = error_TLBuffer_io_in_0_d_valid;
  assign TLBuffer_1_io_out_2_d_bits_opcode = error_TLBuffer_io_in_0_d_bits_opcode;
  assign TLBuffer_1_io_out_2_d_bits_param = error_TLBuffer_io_in_0_d_bits_param;
  assign TLBuffer_1_io_out_2_d_bits_size = error_TLBuffer_io_in_0_d_bits_size;
  assign TLBuffer_1_io_out_2_d_bits_source = error_TLBuffer_io_in_0_d_bits_source;
  assign TLBuffer_1_io_out_2_d_bits_sink = error_TLBuffer_io_in_0_d_bits_sink;
  assign TLBuffer_1_io_out_2_d_bits_data = error_TLBuffer_io_in_0_d_bits_data;
  assign TLBuffer_1_io_out_2_d_bits_error = error_TLBuffer_io_in_0_d_bits_error;
  assign TLBuffer_1_io_out_1_a_ready = TLWidthWidget_io_in_1_a_ready;
  assign TLBuffer_1_io_out_1_d_valid = TLWidthWidget_io_in_1_d_valid;
  assign TLBuffer_1_io_out_1_d_bits_opcode = TLWidthWidget_io_in_1_d_bits_opcode;
  assign TLBuffer_1_io_out_1_d_bits_param = TLWidthWidget_io_in_1_d_bits_param;
  assign TLBuffer_1_io_out_1_d_bits_size = TLWidthWidget_io_in_1_d_bits_size;
  assign TLBuffer_1_io_out_1_d_bits_source = TLWidthWidget_io_in_1_d_bits_source;
  assign TLBuffer_1_io_out_1_d_bits_sink = TLWidthWidget_io_in_1_d_bits_sink;
  assign TLBuffer_1_io_out_1_d_bits_data = TLWidthWidget_io_in_1_d_bits_data;
  assign TLBuffer_1_io_out_1_d_bits_error = TLWidthWidget_io_in_1_d_bits_error;
  assign TLBuffer_1_io_out_0_a_ready = TLWidthWidget_io_in_0_a_ready;
  assign TLBuffer_1_io_out_0_d_valid = TLWidthWidget_io_in_0_d_valid;
  assign TLBuffer_1_io_out_0_d_bits_opcode = TLWidthWidget_io_in_0_d_bits_opcode;
  assign TLBuffer_1_io_out_0_d_bits_param = TLWidthWidget_io_in_0_d_bits_param;
  assign TLBuffer_1_io_out_0_d_bits_size = TLWidthWidget_io_in_0_d_bits_size;
  assign TLBuffer_1_io_out_0_d_bits_source = TLWidthWidget_io_in_0_d_bits_source;
  assign TLBuffer_1_io_out_0_d_bits_sink = TLWidthWidget_io_in_0_d_bits_sink;
  assign TLBuffer_1_io_out_0_d_bits_data = TLWidthWidget_io_in_0_d_bits_data;
  assign TLBuffer_1_io_out_0_d_bits_error = TLWidthWidget_io_in_0_d_bits_error;
  assign TLWidthWidget_clock = clock;
  assign TLWidthWidget_reset = reset;
  assign TLWidthWidget_io_in_1_a_valid = TLBuffer_1_io_out_1_a_valid;
  assign TLWidthWidget_io_in_1_a_bits_opcode = TLBuffer_1_io_out_1_a_bits_opcode;
  assign TLWidthWidget_io_in_1_a_bits_size = TLBuffer_1_io_out_1_a_bits_size;
  assign TLWidthWidget_io_in_1_a_bits_source = TLBuffer_1_io_out_1_a_bits_source;
  assign TLWidthWidget_io_in_1_a_bits_address = TLBuffer_1_io_out_1_a_bits_address;
  assign TLWidthWidget_io_in_1_a_bits_mask = TLBuffer_1_io_out_1_a_bits_mask;
  assign TLWidthWidget_io_in_1_a_bits_data = TLBuffer_1_io_out_1_a_bits_data;
  assign TLWidthWidget_io_in_1_d_ready = TLBuffer_1_io_out_1_d_ready;
  assign TLWidthWidget_io_in_0_a_valid = TLBuffer_1_io_out_0_a_valid;
  assign TLWidthWidget_io_in_0_a_bits_opcode = TLBuffer_1_io_out_0_a_bits_opcode;
  assign TLWidthWidget_io_in_0_a_bits_param = TLBuffer_1_io_out_0_a_bits_param;
  assign TLWidthWidget_io_in_0_a_bits_size = TLBuffer_1_io_out_0_a_bits_size;
  assign TLWidthWidget_io_in_0_a_bits_source = TLBuffer_1_io_out_0_a_bits_source;
  assign TLWidthWidget_io_in_0_a_bits_address = TLBuffer_1_io_out_0_a_bits_address;
  assign TLWidthWidget_io_in_0_a_bits_mask = TLBuffer_1_io_out_0_a_bits_mask;
  assign TLWidthWidget_io_in_0_a_bits_data = TLBuffer_1_io_out_0_a_bits_data;
  assign TLWidthWidget_io_in_0_d_ready = TLBuffer_1_io_out_0_d_ready;
  assign TLWidthWidget_io_out_1_a_ready = TLToAXI4_io_in_0_a_ready;
  assign TLWidthWidget_io_out_1_d_valid = TLToAXI4_io_in_0_d_valid;
  assign TLWidthWidget_io_out_1_d_bits_opcode = TLToAXI4_io_in_0_d_bits_opcode;
  assign TLWidthWidget_io_out_1_d_bits_param = TLToAXI4_io_in_0_d_bits_param;
  assign TLWidthWidget_io_out_1_d_bits_size = TLToAXI4_io_in_0_d_bits_size;
  assign TLWidthWidget_io_out_1_d_bits_source = TLToAXI4_io_in_0_d_bits_source;
  assign TLWidthWidget_io_out_1_d_bits_sink = TLToAXI4_io_in_0_d_bits_sink;
  assign TLWidthWidget_io_out_1_d_bits_data = TLToAXI4_io_in_0_d_bits_data;
  assign TLWidthWidget_io_out_1_d_bits_error = TLToAXI4_io_in_0_d_bits_error;
  assign TLWidthWidget_io_out_0_a_ready = TLAtomicAutomata_io_in_0_a_ready;
  assign TLWidthWidget_io_out_0_d_valid = TLAtomicAutomata_io_in_0_d_valid;
  assign TLWidthWidget_io_out_0_d_bits_opcode = TLAtomicAutomata_io_in_0_d_bits_opcode;
  assign TLWidthWidget_io_out_0_d_bits_param = TLAtomicAutomata_io_in_0_d_bits_param;
  assign TLWidthWidget_io_out_0_d_bits_size = TLAtomicAutomata_io_in_0_d_bits_size;
  assign TLWidthWidget_io_out_0_d_bits_source = TLAtomicAutomata_io_in_0_d_bits_source;
  assign TLWidthWidget_io_out_0_d_bits_sink = TLAtomicAutomata_io_in_0_d_bits_sink;
  assign TLWidthWidget_io_out_0_d_bits_data = TLAtomicAutomata_io_in_0_d_bits_data;
  assign TLWidthWidget_io_out_0_d_bits_error = TLAtomicAutomata_io_in_0_d_bits_error;
  assign TLSplitter_io_in_1_a_valid = TLFIFOFixer_1_io_out_0_a_valid;
  assign TLSplitter_io_in_1_a_bits_opcode = TLFIFOFixer_1_io_out_0_a_bits_opcode;
  assign TLSplitter_io_in_1_a_bits_param = TLFIFOFixer_1_io_out_0_a_bits_param;
  assign TLSplitter_io_in_1_a_bits_size = TLFIFOFixer_1_io_out_0_a_bits_size;
  assign TLSplitter_io_in_1_a_bits_source = TLFIFOFixer_1_io_out_0_a_bits_source;
  assign TLSplitter_io_in_1_a_bits_address = TLFIFOFixer_1_io_out_0_a_bits_address;
  assign TLSplitter_io_in_1_a_bits_mask = TLFIFOFixer_1_io_out_0_a_bits_mask;
  assign TLSplitter_io_in_1_a_bits_data = TLFIFOFixer_1_io_out_0_a_bits_data;
  assign TLSplitter_io_in_1_d_ready = TLFIFOFixer_1_io_out_0_d_ready;
  assign TLSplitter_io_in_0_a_valid = TLFIFOFixer_io_out_0_a_valid;
  assign TLSplitter_io_in_0_a_bits_opcode = TLFIFOFixer_io_out_0_a_bits_opcode;
  assign TLSplitter_io_in_0_a_bits_param = TLFIFOFixer_io_out_0_a_bits_param;
  assign TLSplitter_io_in_0_a_bits_size = TLFIFOFixer_io_out_0_a_bits_size;
  assign TLSplitter_io_in_0_a_bits_source = TLFIFOFixer_io_out_0_a_bits_source;
  assign TLSplitter_io_in_0_a_bits_address = TLFIFOFixer_io_out_0_a_bits_address;
  assign TLSplitter_io_in_0_a_bits_mask = TLFIFOFixer_io_out_0_a_bits_mask;
  assign TLSplitter_io_in_0_a_bits_data = TLFIFOFixer_io_out_0_a_bits_data;
  assign TLSplitter_io_in_0_d_ready = TLFIFOFixer_io_out_0_d_ready;
  assign TLSplitter_io_out_1_a_ready = TLXbar_io_in_1_a_ready;
  assign TLSplitter_io_out_1_d_valid = TLXbar_io_in_1_d_valid;
  assign TLSplitter_io_out_1_d_bits_opcode = TLXbar_io_in_1_d_bits_opcode;
  assign TLSplitter_io_out_1_d_bits_size = TLXbar_io_in_1_d_bits_size;
  assign TLSplitter_io_out_1_d_bits_source = TLXbar_io_in_1_d_bits_source;
  assign TLSplitter_io_out_0_a_ready = TLXbar_io_in_0_a_ready;
  assign TLSplitter_io_out_0_d_valid = TLXbar_io_in_0_d_valid;
  assign TLSplitter_io_out_0_d_bits_opcode = TLXbar_io_in_0_d_bits_opcode;
  assign TLSplitter_io_out_0_d_bits_size = TLXbar_io_in_0_d_bits_size;
  assign TLSplitter_io_out_0_d_bits_source = TLXbar_io_in_0_d_bits_source;
  assign TLSplitter_io_out_0_d_bits_data = TLXbar_io_in_0_d_bits_data;
  assign TLSplitter_io_out_0_d_bits_error = TLXbar_io_in_0_d_bits_error;
  assign TLFIFOFixer_io_in_0_a_valid = TLBuffer_4_io_out_0_a_valid;
  assign TLFIFOFixer_io_in_0_a_bits_opcode = TLBuffer_4_io_out_0_a_bits_opcode;
  assign TLFIFOFixer_io_in_0_a_bits_param = TLBuffer_4_io_out_0_a_bits_param;
  assign TLFIFOFixer_io_in_0_a_bits_size = TLBuffer_4_io_out_0_a_bits_size;
  assign TLFIFOFixer_io_in_0_a_bits_source = TLBuffer_4_io_out_0_a_bits_source;
  assign TLFIFOFixer_io_in_0_a_bits_address = TLBuffer_4_io_out_0_a_bits_address;
  assign TLFIFOFixer_io_in_0_a_bits_mask = TLBuffer_4_io_out_0_a_bits_mask;
  assign TLFIFOFixer_io_in_0_a_bits_data = TLBuffer_4_io_out_0_a_bits_data;
  assign TLFIFOFixer_io_in_0_d_ready = TLBuffer_4_io_out_0_d_ready;
  assign TLFIFOFixer_io_out_0_a_ready = TLSplitter_io_in_0_a_ready;
  assign TLFIFOFixer_io_out_0_d_valid = TLSplitter_io_in_0_d_valid;
  assign TLFIFOFixer_io_out_0_d_bits_opcode = TLSplitter_io_in_0_d_bits_opcode;
  assign TLFIFOFixer_io_out_0_d_bits_size = TLSplitter_io_in_0_d_bits_size;
  assign TLFIFOFixer_io_out_0_d_bits_source = TLSplitter_io_in_0_d_bits_source;
  assign TLFIFOFixer_io_out_0_d_bits_data = TLSplitter_io_in_0_d_bits_data;
  assign TLFIFOFixer_io_out_0_d_bits_error = TLSplitter_io_in_0_d_bits_error;
  assign TLFIFOFixer_1_clock = clock;
  assign TLFIFOFixer_1_reset = reset;
  assign TLFIFOFixer_1_io_in_0_a_valid = TLBuffer_5_io_out_0_a_valid;
  assign TLFIFOFixer_1_io_in_0_a_bits_opcode = TLBuffer_5_io_out_0_a_bits_opcode;
  assign TLFIFOFixer_1_io_in_0_a_bits_param = TLBuffer_5_io_out_0_a_bits_param;
  assign TLFIFOFixer_1_io_in_0_a_bits_size = TLBuffer_5_io_out_0_a_bits_size;
  assign TLFIFOFixer_1_io_in_0_a_bits_source = TLBuffer_5_io_out_0_a_bits_source;
  assign TLFIFOFixer_1_io_in_0_a_bits_address = TLBuffer_5_io_out_0_a_bits_address;
  assign TLFIFOFixer_1_io_in_0_a_bits_mask = TLBuffer_5_io_out_0_a_bits_mask;
  assign TLFIFOFixer_1_io_in_0_a_bits_data = TLBuffer_5_io_out_0_a_bits_data;
  assign TLFIFOFixer_1_io_in_0_d_ready = TLBuffer_5_io_out_0_d_ready;
  assign TLFIFOFixer_1_io_out_0_a_ready = TLSplitter_io_in_1_a_ready;
  assign TLFIFOFixer_1_io_out_0_d_valid = TLSplitter_io_in_1_d_valid;
  assign TLFIFOFixer_1_io_out_0_d_bits_opcode = TLSplitter_io_in_1_d_bits_opcode;
  assign TLFIFOFixer_1_io_out_0_d_bits_size = TLSplitter_io_in_1_d_bits_size;
  assign TLFIFOFixer_1_io_out_0_d_bits_source = TLSplitter_io_in_1_d_bits_source;
  assign TLXbar_1_clock = clock;
  assign TLXbar_1_reset = reset;
  assign TLXbar_1_io_in_0_a_valid = TLBuffer_2_io_out_0_a_valid;
  assign TLXbar_1_io_in_0_a_bits_opcode = TLBuffer_2_io_out_0_a_bits_opcode;
  assign TLXbar_1_io_in_0_a_bits_param = TLBuffer_2_io_out_0_a_bits_param;
  assign TLXbar_1_io_in_0_a_bits_size = TLBuffer_2_io_out_0_a_bits_size;
  assign TLXbar_1_io_in_0_a_bits_source = TLBuffer_2_io_out_0_a_bits_source;
  assign TLXbar_1_io_in_0_a_bits_address = TLBuffer_2_io_out_0_a_bits_address;
  assign TLXbar_1_io_in_0_a_bits_mask = TLBuffer_2_io_out_0_a_bits_mask;
  assign TLXbar_1_io_in_0_a_bits_data = TLBuffer_2_io_out_0_a_bits_data;
  assign TLXbar_1_io_in_0_d_ready = TLBuffer_2_io_out_0_d_ready;
  assign TLXbar_1_io_out_4_a_ready = TLBuffer_3_io_in_4_a_ready;
  assign TLXbar_1_io_out_4_d_valid = TLBuffer_3_io_in_4_d_valid;
  assign TLXbar_1_io_out_4_d_bits_opcode = TLBuffer_3_io_in_4_d_bits_opcode;
  assign TLXbar_1_io_out_4_d_bits_param = TLBuffer_3_io_in_4_d_bits_param;
  assign TLXbar_1_io_out_4_d_bits_size = TLBuffer_3_io_in_4_d_bits_size;
  assign TLXbar_1_io_out_4_d_bits_source = TLBuffer_3_io_in_4_d_bits_source;
  assign TLXbar_1_io_out_4_d_bits_sink = TLBuffer_3_io_in_4_d_bits_sink;
  assign TLXbar_1_io_out_4_d_bits_data = TLBuffer_3_io_in_4_d_bits_data;
  assign TLXbar_1_io_out_4_d_bits_error = TLBuffer_3_io_in_4_d_bits_error;
  assign TLXbar_1_io_out_3_a_ready = TLBuffer_3_io_in_3_a_ready;
  assign TLXbar_1_io_out_3_d_valid = TLBuffer_3_io_in_3_d_valid;
  assign TLXbar_1_io_out_3_d_bits_opcode = TLBuffer_3_io_in_3_d_bits_opcode;
  assign TLXbar_1_io_out_3_d_bits_param = TLBuffer_3_io_in_3_d_bits_param;
  assign TLXbar_1_io_out_3_d_bits_size = TLBuffer_3_io_in_3_d_bits_size;
  assign TLXbar_1_io_out_3_d_bits_source = TLBuffer_3_io_in_3_d_bits_source;
  assign TLXbar_1_io_out_3_d_bits_sink = TLBuffer_3_io_in_3_d_bits_sink;
  assign TLXbar_1_io_out_3_d_bits_data = TLBuffer_3_io_in_3_d_bits_data;
  assign TLXbar_1_io_out_3_d_bits_error = TLBuffer_3_io_in_3_d_bits_error;
  assign TLXbar_1_io_out_2_a_ready = TLBuffer_3_io_in_2_a_ready;
  assign TLXbar_1_io_out_2_d_valid = TLBuffer_3_io_in_2_d_valid;
  assign TLXbar_1_io_out_2_d_bits_opcode = TLBuffer_3_io_in_2_d_bits_opcode;
  assign TLXbar_1_io_out_2_d_bits_param = TLBuffer_3_io_in_2_d_bits_param;
  assign TLXbar_1_io_out_2_d_bits_size = TLBuffer_3_io_in_2_d_bits_size;
  assign TLXbar_1_io_out_2_d_bits_source = TLBuffer_3_io_in_2_d_bits_source;
  assign TLXbar_1_io_out_2_d_bits_sink = TLBuffer_3_io_in_2_d_bits_sink;
  assign TLXbar_1_io_out_2_d_bits_data = TLBuffer_3_io_in_2_d_bits_data;
  assign TLXbar_1_io_out_2_d_bits_error = TLBuffer_3_io_in_2_d_bits_error;
  assign TLXbar_1_io_out_1_a_ready = TLBuffer_3_io_in_1_a_ready;
  assign TLXbar_1_io_out_1_d_valid = TLBuffer_3_io_in_1_d_valid;
  assign TLXbar_1_io_out_1_d_bits_opcode = TLBuffer_3_io_in_1_d_bits_opcode;
  assign TLXbar_1_io_out_1_d_bits_param = TLBuffer_3_io_in_1_d_bits_param;
  assign TLXbar_1_io_out_1_d_bits_size = TLBuffer_3_io_in_1_d_bits_size;
  assign TLXbar_1_io_out_1_d_bits_source = TLBuffer_3_io_in_1_d_bits_source;
  assign TLXbar_1_io_out_1_d_bits_sink = TLBuffer_3_io_in_1_d_bits_sink;
  assign TLXbar_1_io_out_1_d_bits_data = TLBuffer_3_io_in_1_d_bits_data;
  assign TLXbar_1_io_out_1_d_bits_error = TLBuffer_3_io_in_1_d_bits_error;
  assign TLXbar_1_io_out_0_a_ready = TLBuffer_3_io_in_0_a_ready;
  assign TLXbar_1_io_out_0_d_valid = TLBuffer_3_io_in_0_d_valid;
  assign TLXbar_1_io_out_0_d_bits_opcode = TLBuffer_3_io_in_0_d_bits_opcode;
  assign TLXbar_1_io_out_0_d_bits_param = TLBuffer_3_io_in_0_d_bits_param;
  assign TLXbar_1_io_out_0_d_bits_size = TLBuffer_3_io_in_0_d_bits_size;
  assign TLXbar_1_io_out_0_d_bits_source = TLBuffer_3_io_in_0_d_bits_source;
  assign TLXbar_1_io_out_0_d_bits_sink = TLBuffer_3_io_in_0_d_bits_sink;
  assign TLXbar_1_io_out_0_d_bits_data = TLBuffer_3_io_in_0_d_bits_data;
  assign TLXbar_1_io_out_0_d_bits_error = TLBuffer_3_io_in_0_d_bits_error;
  assign TLBuffer_2_clock = clock;
  assign TLBuffer_2_reset = reset;
  assign TLBuffer_2_io_in_0_a_valid = TLAtomicAutomata_io_out_0_a_valid;
  assign TLBuffer_2_io_in_0_a_bits_opcode = TLAtomicAutomata_io_out_0_a_bits_opcode;
  assign TLBuffer_2_io_in_0_a_bits_param = TLAtomicAutomata_io_out_0_a_bits_param;
  assign TLBuffer_2_io_in_0_a_bits_size = TLAtomicAutomata_io_out_0_a_bits_size;
  assign TLBuffer_2_io_in_0_a_bits_source = TLAtomicAutomata_io_out_0_a_bits_source;
  assign TLBuffer_2_io_in_0_a_bits_address = TLAtomicAutomata_io_out_0_a_bits_address;
  assign TLBuffer_2_io_in_0_a_bits_mask = TLAtomicAutomata_io_out_0_a_bits_mask;
  assign TLBuffer_2_io_in_0_a_bits_data = TLAtomicAutomata_io_out_0_a_bits_data;
  assign TLBuffer_2_io_in_0_d_ready = TLAtomicAutomata_io_out_0_d_ready;
  assign TLBuffer_2_io_out_0_a_ready = TLXbar_1_io_in_0_a_ready;
  assign TLBuffer_2_io_out_0_d_valid = TLXbar_1_io_in_0_d_valid;
  assign TLBuffer_2_io_out_0_d_bits_opcode = TLXbar_1_io_in_0_d_bits_opcode;
  assign TLBuffer_2_io_out_0_d_bits_param = TLXbar_1_io_in_0_d_bits_param;
  assign TLBuffer_2_io_out_0_d_bits_size = TLXbar_1_io_in_0_d_bits_size;
  assign TLBuffer_2_io_out_0_d_bits_source = TLXbar_1_io_in_0_d_bits_source;
  assign TLBuffer_2_io_out_0_d_bits_sink = TLXbar_1_io_in_0_d_bits_sink;
  assign TLBuffer_2_io_out_0_d_bits_data = TLXbar_1_io_in_0_d_bits_data;
  assign TLBuffer_2_io_out_0_d_bits_error = TLXbar_1_io_in_0_d_bits_error;
  assign TLBuffer_3_io_in_4_a_valid = TLXbar_1_io_out_4_a_valid;
  assign TLBuffer_3_io_in_4_a_bits_opcode = TLXbar_1_io_out_4_a_bits_opcode;
  assign TLBuffer_3_io_in_4_a_bits_param = TLXbar_1_io_out_4_a_bits_param;
  assign TLBuffer_3_io_in_4_a_bits_size = TLXbar_1_io_out_4_a_bits_size;
  assign TLBuffer_3_io_in_4_a_bits_source = TLXbar_1_io_out_4_a_bits_source;
  assign TLBuffer_3_io_in_4_a_bits_address = TLXbar_1_io_out_4_a_bits_address;
  assign TLBuffer_3_io_in_4_a_bits_mask = TLXbar_1_io_out_4_a_bits_mask;
  assign TLBuffer_3_io_in_4_a_bits_data = TLXbar_1_io_out_4_a_bits_data;
  assign TLBuffer_3_io_in_4_d_ready = TLXbar_1_io_out_4_d_ready;
  assign TLBuffer_3_io_in_3_a_valid = TLXbar_1_io_out_3_a_valid;
  assign TLBuffer_3_io_in_3_a_bits_opcode = TLXbar_1_io_out_3_a_bits_opcode;
  assign TLBuffer_3_io_in_3_a_bits_size = TLXbar_1_io_out_3_a_bits_size;
  assign TLBuffer_3_io_in_3_a_bits_source = TLXbar_1_io_out_3_a_bits_source;
  assign TLBuffer_3_io_in_3_a_bits_address = TLXbar_1_io_out_3_a_bits_address;
  assign TLBuffer_3_io_in_3_a_bits_mask = TLXbar_1_io_out_3_a_bits_mask;
  assign TLBuffer_3_io_in_3_d_ready = TLXbar_1_io_out_3_d_ready;
  assign TLBuffer_3_io_in_2_a_valid = TLXbar_1_io_out_2_a_valid;
  assign TLBuffer_3_io_in_2_a_bits_opcode = TLXbar_1_io_out_2_a_bits_opcode;
  assign TLBuffer_3_io_in_2_a_bits_size = TLXbar_1_io_out_2_a_bits_size;
  assign TLBuffer_3_io_in_2_a_bits_source = TLXbar_1_io_out_2_a_bits_source;
  assign TLBuffer_3_io_in_2_a_bits_address = TLXbar_1_io_out_2_a_bits_address;
  assign TLBuffer_3_io_in_2_a_bits_mask = TLXbar_1_io_out_2_a_bits_mask;
  assign TLBuffer_3_io_in_2_a_bits_data = TLXbar_1_io_out_2_a_bits_data;
  assign TLBuffer_3_io_in_2_d_ready = TLXbar_1_io_out_2_d_ready;
  assign TLBuffer_3_io_in_1_a_valid = TLXbar_1_io_out_1_a_valid;
  assign TLBuffer_3_io_in_1_a_bits_opcode = TLXbar_1_io_out_1_a_bits_opcode;
  assign TLBuffer_3_io_in_1_a_bits_size = TLXbar_1_io_out_1_a_bits_size;
  assign TLBuffer_3_io_in_1_a_bits_source = TLXbar_1_io_out_1_a_bits_source;
  assign TLBuffer_3_io_in_1_a_bits_address = TLXbar_1_io_out_1_a_bits_address;
  assign TLBuffer_3_io_in_1_a_bits_mask = TLXbar_1_io_out_1_a_bits_mask;
  assign TLBuffer_3_io_in_1_a_bits_data = TLXbar_1_io_out_1_a_bits_data;
  assign TLBuffer_3_io_in_1_d_ready = TLXbar_1_io_out_1_d_ready;
  assign TLBuffer_3_io_in_0_a_valid = TLXbar_1_io_out_0_a_valid;
  assign TLBuffer_3_io_in_0_a_bits_opcode = TLXbar_1_io_out_0_a_bits_opcode;
  assign TLBuffer_3_io_in_0_a_bits_size = TLXbar_1_io_out_0_a_bits_size;
  assign TLBuffer_3_io_in_0_a_bits_source = TLXbar_1_io_out_0_a_bits_source;
  assign TLBuffer_3_io_in_0_a_bits_address = TLXbar_1_io_out_0_a_bits_address;
  assign TLBuffer_3_io_in_0_a_bits_mask = TLXbar_1_io_out_0_a_bits_mask;
  assign TLBuffer_3_io_in_0_a_bits_data = TLXbar_1_io_out_0_a_bits_data;
  assign TLBuffer_3_io_in_0_d_ready = TLXbar_1_io_out_0_d_ready;
  assign TLBuffer_3_io_out_4_a_ready = tile_io_slave_0_a_ready;
  assign TLBuffer_3_io_out_4_d_valid = tile_io_slave_0_d_valid;
  assign TLBuffer_3_io_out_4_d_bits_opcode = tile_io_slave_0_d_bits_opcode;
  assign TLBuffer_3_io_out_4_d_bits_param = tile_io_slave_0_d_bits_param;
  assign TLBuffer_3_io_out_4_d_bits_size = tile_io_slave_0_d_bits_size;
  assign TLBuffer_3_io_out_4_d_bits_source = tile_io_slave_0_d_bits_source;
  assign TLBuffer_3_io_out_4_d_bits_sink = tile_io_slave_0_d_bits_sink;
  assign TLBuffer_3_io_out_4_d_bits_data = tile_io_slave_0_d_bits_data;
  assign TLBuffer_3_io_out_4_d_bits_error = tile_io_slave_0_d_bits_error;
  assign TLBuffer_3_io_out_3_a_ready = TLFragmenter_1_io_in_3_a_ready;
  assign TLBuffer_3_io_out_3_d_valid = TLFragmenter_1_io_in_3_d_valid;
  assign TLBuffer_3_io_out_3_d_bits_opcode = TLFragmenter_1_io_in_3_d_bits_opcode;
  assign TLBuffer_3_io_out_3_d_bits_param = TLFragmenter_1_io_in_3_d_bits_param;
  assign TLBuffer_3_io_out_3_d_bits_size = TLFragmenter_1_io_in_3_d_bits_size;
  assign TLBuffer_3_io_out_3_d_bits_source = TLFragmenter_1_io_in_3_d_bits_source;
  assign TLBuffer_3_io_out_3_d_bits_sink = TLFragmenter_1_io_in_3_d_bits_sink;
  assign TLBuffer_3_io_out_3_d_bits_data = TLFragmenter_1_io_in_3_d_bits_data;
  assign TLBuffer_3_io_out_3_d_bits_error = TLFragmenter_1_io_in_3_d_bits_error;
  assign TLBuffer_3_io_out_2_a_ready = TLFragmenter_1_io_in_2_a_ready;
  assign TLBuffer_3_io_out_2_d_valid = TLFragmenter_1_io_in_2_d_valid;
  assign TLBuffer_3_io_out_2_d_bits_opcode = TLFragmenter_1_io_in_2_d_bits_opcode;
  assign TLBuffer_3_io_out_2_d_bits_param = TLFragmenter_1_io_in_2_d_bits_param;
  assign TLBuffer_3_io_out_2_d_bits_size = TLFragmenter_1_io_in_2_d_bits_size;
  assign TLBuffer_3_io_out_2_d_bits_source = TLFragmenter_1_io_in_2_d_bits_source;
  assign TLBuffer_3_io_out_2_d_bits_sink = TLFragmenter_1_io_in_2_d_bits_sink;
  assign TLBuffer_3_io_out_2_d_bits_data = TLFragmenter_1_io_in_2_d_bits_data;
  assign TLBuffer_3_io_out_2_d_bits_error = TLFragmenter_1_io_in_2_d_bits_error;
  assign TLBuffer_3_io_out_1_a_ready = TLFragmenter_1_io_in_1_a_ready;
  assign TLBuffer_3_io_out_1_d_valid = TLFragmenter_1_io_in_1_d_valid;
  assign TLBuffer_3_io_out_1_d_bits_opcode = TLFragmenter_1_io_in_1_d_bits_opcode;
  assign TLBuffer_3_io_out_1_d_bits_param = TLFragmenter_1_io_in_1_d_bits_param;
  assign TLBuffer_3_io_out_1_d_bits_size = TLFragmenter_1_io_in_1_d_bits_size;
  assign TLBuffer_3_io_out_1_d_bits_source = TLFragmenter_1_io_in_1_d_bits_source;
  assign TLBuffer_3_io_out_1_d_bits_sink = TLFragmenter_1_io_in_1_d_bits_sink;
  assign TLBuffer_3_io_out_1_d_bits_data = TLFragmenter_1_io_in_1_d_bits_data;
  assign TLBuffer_3_io_out_1_d_bits_error = TLFragmenter_1_io_in_1_d_bits_error;
  assign TLBuffer_3_io_out_0_a_ready = TLFragmenter_1_io_in_0_a_ready;
  assign TLBuffer_3_io_out_0_d_valid = TLFragmenter_1_io_in_0_d_valid;
  assign TLBuffer_3_io_out_0_d_bits_opcode = TLFragmenter_1_io_in_0_d_bits_opcode;
  assign TLBuffer_3_io_out_0_d_bits_param = TLFragmenter_1_io_in_0_d_bits_param;
  assign TLBuffer_3_io_out_0_d_bits_size = TLFragmenter_1_io_in_0_d_bits_size;
  assign TLBuffer_3_io_out_0_d_bits_source = TLFragmenter_1_io_in_0_d_bits_source;
  assign TLBuffer_3_io_out_0_d_bits_sink = TLFragmenter_1_io_in_0_d_bits_sink;
  assign TLBuffer_3_io_out_0_d_bits_data = TLFragmenter_1_io_in_0_d_bits_data;
  assign TLBuffer_3_io_out_0_d_bits_error = TLFragmenter_1_io_in_0_d_bits_error;
  assign TLFragmenter_1_clock = clock;
  assign TLFragmenter_1_reset = reset;
  assign TLFragmenter_1_io_in_3_a_valid = TLBuffer_3_io_out_3_a_valid;
  assign TLFragmenter_1_io_in_3_a_bits_opcode = TLBuffer_3_io_out_3_a_bits_opcode;
  assign TLFragmenter_1_io_in_3_a_bits_size = TLBuffer_3_io_out_3_a_bits_size;
  assign TLFragmenter_1_io_in_3_a_bits_source = TLBuffer_3_io_out_3_a_bits_source;
  assign TLFragmenter_1_io_in_3_a_bits_address = TLBuffer_3_io_out_3_a_bits_address;
  assign TLFragmenter_1_io_in_3_a_bits_mask = TLBuffer_3_io_out_3_a_bits_mask;
  assign TLFragmenter_1_io_in_3_d_ready = TLBuffer_3_io_out_3_d_ready;
  assign TLFragmenter_1_io_in_2_a_valid = TLBuffer_3_io_out_2_a_valid;
  assign TLFragmenter_1_io_in_2_a_bits_opcode = TLBuffer_3_io_out_2_a_bits_opcode;
  assign TLFragmenter_1_io_in_2_a_bits_size = TLBuffer_3_io_out_2_a_bits_size;
  assign TLFragmenter_1_io_in_2_a_bits_source = TLBuffer_3_io_out_2_a_bits_source;
  assign TLFragmenter_1_io_in_2_a_bits_address = TLBuffer_3_io_out_2_a_bits_address;
  assign TLFragmenter_1_io_in_2_a_bits_mask = TLBuffer_3_io_out_2_a_bits_mask;
  assign TLFragmenter_1_io_in_2_a_bits_data = TLBuffer_3_io_out_2_a_bits_data;
  assign TLFragmenter_1_io_in_2_d_ready = TLBuffer_3_io_out_2_d_ready;
  assign TLFragmenter_1_io_in_1_a_valid = TLBuffer_3_io_out_1_a_valid;
  assign TLFragmenter_1_io_in_1_a_bits_opcode = TLBuffer_3_io_out_1_a_bits_opcode;
  assign TLFragmenter_1_io_in_1_a_bits_size = TLBuffer_3_io_out_1_a_bits_size;
  assign TLFragmenter_1_io_in_1_a_bits_source = TLBuffer_3_io_out_1_a_bits_source;
  assign TLFragmenter_1_io_in_1_a_bits_address = TLBuffer_3_io_out_1_a_bits_address;
  assign TLFragmenter_1_io_in_1_a_bits_mask = TLBuffer_3_io_out_1_a_bits_mask;
  assign TLFragmenter_1_io_in_1_a_bits_data = TLBuffer_3_io_out_1_a_bits_data;
  assign TLFragmenter_1_io_in_1_d_ready = TLBuffer_3_io_out_1_d_ready;
  assign TLFragmenter_1_io_in_0_a_valid = TLBuffer_3_io_out_0_a_valid;
  assign TLFragmenter_1_io_in_0_a_bits_opcode = TLBuffer_3_io_out_0_a_bits_opcode;
  assign TLFragmenter_1_io_in_0_a_bits_size = TLBuffer_3_io_out_0_a_bits_size;
  assign TLFragmenter_1_io_in_0_a_bits_source = TLBuffer_3_io_out_0_a_bits_source;
  assign TLFragmenter_1_io_in_0_a_bits_address = TLBuffer_3_io_out_0_a_bits_address;
  assign TLFragmenter_1_io_in_0_a_bits_mask = TLBuffer_3_io_out_0_a_bits_mask;
  assign TLFragmenter_1_io_in_0_a_bits_data = TLBuffer_3_io_out_0_a_bits_data;
  assign TLFragmenter_1_io_in_0_d_ready = TLBuffer_3_io_out_0_d_ready;
  assign TLFragmenter_1_io_out_3_a_ready = bootrom_io_in_0_a_ready;
  assign TLFragmenter_1_io_out_3_d_valid = bootrom_io_in_0_d_valid;
  assign TLFragmenter_1_io_out_3_d_bits_opcode = bootrom_io_in_0_d_bits_opcode;
  assign TLFragmenter_1_io_out_3_d_bits_param = bootrom_io_in_0_d_bits_param;
  assign TLFragmenter_1_io_out_3_d_bits_size = bootrom_io_in_0_d_bits_size;
  assign TLFragmenter_1_io_out_3_d_bits_source = bootrom_io_in_0_d_bits_source;
  assign TLFragmenter_1_io_out_3_d_bits_sink = bootrom_io_in_0_d_bits_sink;
  assign TLFragmenter_1_io_out_3_d_bits_data = bootrom_io_in_0_d_bits_data;
  assign TLFragmenter_1_io_out_3_d_bits_error = bootrom_io_in_0_d_bits_error;
  assign TLFragmenter_1_io_out_2_a_ready = debug_1_io_in_0_a_ready;
  assign TLFragmenter_1_io_out_2_d_valid = debug_1_io_in_0_d_valid;
  assign TLFragmenter_1_io_out_2_d_bits_opcode = debug_1_io_in_0_d_bits_opcode;
  assign TLFragmenter_1_io_out_2_d_bits_param = debug_1_io_in_0_d_bits_param;
  assign TLFragmenter_1_io_out_2_d_bits_size = debug_1_io_in_0_d_bits_size;
  assign TLFragmenter_1_io_out_2_d_bits_source = debug_1_io_in_0_d_bits_source;
  assign TLFragmenter_1_io_out_2_d_bits_sink = debug_1_io_in_0_d_bits_sink;
  assign TLFragmenter_1_io_out_2_d_bits_data = debug_1_io_in_0_d_bits_data;
  assign TLFragmenter_1_io_out_2_d_bits_error = debug_1_io_in_0_d_bits_error;
  assign TLFragmenter_1_io_out_1_a_ready = clint_io_in_0_a_ready;
  assign TLFragmenter_1_io_out_1_d_valid = clint_io_in_0_d_valid;
  assign TLFragmenter_1_io_out_1_d_bits_opcode = clint_io_in_0_d_bits_opcode;
  assign TLFragmenter_1_io_out_1_d_bits_param = clint_io_in_0_d_bits_param;
  assign TLFragmenter_1_io_out_1_d_bits_size = clint_io_in_0_d_bits_size;
  assign TLFragmenter_1_io_out_1_d_bits_source = clint_io_in_0_d_bits_source;
  assign TLFragmenter_1_io_out_1_d_bits_sink = clint_io_in_0_d_bits_sink;
  assign TLFragmenter_1_io_out_1_d_bits_data = clint_io_in_0_d_bits_data;
  assign TLFragmenter_1_io_out_1_d_bits_error = clint_io_in_0_d_bits_error;
  assign TLFragmenter_1_io_out_0_a_ready = plic_io_tl_in_0_a_ready;
  assign TLFragmenter_1_io_out_0_d_valid = plic_io_tl_in_0_d_valid;
  assign TLFragmenter_1_io_out_0_d_bits_opcode = plic_io_tl_in_0_d_bits_opcode;
  assign TLFragmenter_1_io_out_0_d_bits_param = plic_io_tl_in_0_d_bits_param;
  assign TLFragmenter_1_io_out_0_d_bits_size = plic_io_tl_in_0_d_bits_size;
  assign TLFragmenter_1_io_out_0_d_bits_source = plic_io_tl_in_0_d_bits_source;
  assign TLFragmenter_1_io_out_0_d_bits_sink = plic_io_tl_in_0_d_bits_sink;
  assign TLFragmenter_1_io_out_0_d_bits_data = plic_io_tl_in_0_d_bits_data;
  assign TLFragmenter_1_io_out_0_d_bits_error = plic_io_tl_in_0_d_bits_error;
  assign TLAtomicAutomata_clock = clock;
  assign TLAtomicAutomata_reset = reset;
  assign TLAtomicAutomata_io_in_0_a_valid = TLWidthWidget_io_out_0_a_valid;
  assign TLAtomicAutomata_io_in_0_a_bits_opcode = TLWidthWidget_io_out_0_a_bits_opcode;
  assign TLAtomicAutomata_io_in_0_a_bits_param = TLWidthWidget_io_out_0_a_bits_param;
  assign TLAtomicAutomata_io_in_0_a_bits_size = TLWidthWidget_io_out_0_a_bits_size;
  assign TLAtomicAutomata_io_in_0_a_bits_source = TLWidthWidget_io_out_0_a_bits_source;
  assign TLAtomicAutomata_io_in_0_a_bits_address = TLWidthWidget_io_out_0_a_bits_address;
  assign TLAtomicAutomata_io_in_0_a_bits_mask = TLWidthWidget_io_out_0_a_bits_mask;
  assign TLAtomicAutomata_io_in_0_a_bits_data = TLWidthWidget_io_out_0_a_bits_data;
  assign TLAtomicAutomata_io_in_0_d_ready = TLWidthWidget_io_out_0_d_ready;
  assign TLAtomicAutomata_io_out_0_a_ready = TLBuffer_2_io_in_0_a_ready;
  assign TLAtomicAutomata_io_out_0_d_valid = TLBuffer_2_io_in_0_d_valid;
  assign TLAtomicAutomata_io_out_0_d_bits_opcode = TLBuffer_2_io_in_0_d_bits_opcode;
  assign TLAtomicAutomata_io_out_0_d_bits_param = TLBuffer_2_io_in_0_d_bits_param;
  assign TLAtomicAutomata_io_out_0_d_bits_size = TLBuffer_2_io_in_0_d_bits_size;
  assign TLAtomicAutomata_io_out_0_d_bits_source = TLBuffer_2_io_in_0_d_bits_source;
  assign TLAtomicAutomata_io_out_0_d_bits_sink = TLBuffer_2_io_in_0_d_bits_sink;
  assign TLAtomicAutomata_io_out_0_d_bits_data = TLBuffer_2_io_in_0_d_bits_data;
  assign TLAtomicAutomata_io_out_0_d_bits_error = TLBuffer_2_io_in_0_d_bits_error;
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io_tl_in_0_a_valid = TLFragmenter_1_io_out_0_a_valid;
  assign plic_io_tl_in_0_a_bits_opcode = TLFragmenter_1_io_out_0_a_bits_opcode;
  assign plic_io_tl_in_0_a_bits_size = TLFragmenter_1_io_out_0_a_bits_size;
  assign plic_io_tl_in_0_a_bits_source = TLFragmenter_1_io_out_0_a_bits_source;
  assign plic_io_tl_in_0_a_bits_address = TLFragmenter_1_io_out_0_a_bits_address;
  assign plic_io_tl_in_0_a_bits_mask = TLFragmenter_1_io_out_0_a_bits_mask;
  assign plic_io_tl_in_0_a_bits_data = TLFragmenter_1_io_out_0_a_bits_data;
  assign plic_io_tl_in_0_d_ready = TLFragmenter_1_io_out_0_d_ready;
  assign plic_io_devices_0_0 = IntXbar_io_out_0_0;
  assign plic_io_devices_0_1 = IntXbar_io_out_0_1;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_rtcTick = _T_158;
  assign clint_io_in_0_a_valid = TLFragmenter_1_io_out_1_a_valid;
  assign clint_io_in_0_a_bits_opcode = TLFragmenter_1_io_out_1_a_bits_opcode;
  assign clint_io_in_0_a_bits_size = TLFragmenter_1_io_out_1_a_bits_size;
  assign clint_io_in_0_a_bits_source = TLFragmenter_1_io_out_1_a_bits_source;
  assign clint_io_in_0_a_bits_address = TLFragmenter_1_io_out_1_a_bits_address;
  assign clint_io_in_0_a_bits_mask = TLFragmenter_1_io_out_1_a_bits_mask;
  assign clint_io_in_0_a_bits_data = TLFragmenter_1_io_out_1_a_bits_data;
  assign clint_io_in_0_d_ready = TLFragmenter_1_io_out_1_d_ready;
  assign debug_1_clock = clock;
  assign debug_1_reset = reset;
  assign debug_1_io_in_0_a_valid = TLFragmenter_1_io_out_2_a_valid;
  assign debug_1_io_in_0_a_bits_opcode = TLFragmenter_1_io_out_2_a_bits_opcode;
  assign debug_1_io_in_0_a_bits_size = TLFragmenter_1_io_out_2_a_bits_size;
  assign debug_1_io_in_0_a_bits_source = TLFragmenter_1_io_out_2_a_bits_source;
  assign debug_1_io_in_0_a_bits_address = TLFragmenter_1_io_out_2_a_bits_address;
  assign debug_1_io_in_0_a_bits_mask = TLFragmenter_1_io_out_2_a_bits_mask;
  assign debug_1_io_in_0_a_bits_data = TLFragmenter_1_io_out_2_a_bits_data;
  assign debug_1_io_in_0_d_ready = TLFragmenter_1_io_out_2_d_ready;
  assign debug_1_io_ctrl_debugUnavail_0 = 1'h0;
  assign debug_1_io_dmi_dmi_req_valid = debug_clockeddmi_dmi_req_valid;
  assign debug_1_io_dmi_dmi_req_bits_addr = debug_clockeddmi_dmi_req_bits_addr;
  assign debug_1_io_dmi_dmi_req_bits_data = debug_clockeddmi_dmi_req_bits_data;
  assign debug_1_io_dmi_dmi_req_bits_op = debug_clockeddmi_dmi_req_bits_op;
  assign debug_1_io_dmi_dmi_resp_ready = debug_clockeddmi_dmi_resp_ready;
  assign debug_1_io_dmi_dmiClock = debug_clockeddmi_dmiClock;
  assign debug_1_io_dmi_dmiReset = debug_clockeddmi_dmiReset;
  assign tile_clock = clock;
  assign tile_reset = reset;
  assign tile_io_master_0_a_ready = TLBuffer_4_io_in_0_a_ready;
  assign tile_io_master_0_d_valid = TLBuffer_4_io_in_0_d_valid;
  assign tile_io_master_0_d_bits_opcode = TLBuffer_4_io_in_0_d_bits_opcode;
  assign tile_io_master_0_d_bits_size = TLBuffer_4_io_in_0_d_bits_size;
  assign tile_io_master_0_d_bits_source = TLBuffer_4_io_in_0_d_bits_source;
  assign tile_io_master_0_d_bits_data = TLBuffer_4_io_in_0_d_bits_data;
  assign tile_io_master_0_d_bits_error = TLBuffer_4_io_in_0_d_bits_error;
  assign tile_io_slave_0_a_valid = TLBuffer_3_io_out_4_a_valid;
  assign tile_io_slave_0_a_bits_opcode = TLBuffer_3_io_out_4_a_bits_opcode;
  assign tile_io_slave_0_a_bits_param = TLBuffer_3_io_out_4_a_bits_param;
  assign tile_io_slave_0_a_bits_size = TLBuffer_3_io_out_4_a_bits_size;
  assign tile_io_slave_0_a_bits_source = TLBuffer_3_io_out_4_a_bits_source;
  assign tile_io_slave_0_a_bits_address = TLBuffer_3_io_out_4_a_bits_address;
  assign tile_io_slave_0_a_bits_mask = TLBuffer_3_io_out_4_a_bits_mask;
  assign tile_io_slave_0_a_bits_data = TLBuffer_3_io_out_4_a_bits_data;
  assign tile_io_slave_0_d_ready = TLBuffer_3_io_out_4_d_ready;
  assign tile_io_asyncInterrupts_0_0 = IntXbar_1_io_out_0_0;
  assign tile_io_periphInterrupts_0_0 = IntXbar_2_io_out_0_0;
  assign tile_io_periphInterrupts_0_1 = IntXbar_2_io_out_0_1;
  assign tile_io_periphInterrupts_0_2 = IntXbar_2_io_out_0_2;
  assign tile_io_hartid = 1'h0;
  assign tile_io_resetVector = 32'h10040;
  assign TLBuffer_4_clock = clock;
  assign TLBuffer_4_reset = reset;
  assign TLBuffer_4_io_in_0_a_valid = tile_io_master_0_a_valid;
  assign TLBuffer_4_io_in_0_a_bits_opcode = tile_io_master_0_a_bits_opcode;
  assign TLBuffer_4_io_in_0_a_bits_param = tile_io_master_0_a_bits_param;
  assign TLBuffer_4_io_in_0_a_bits_size = tile_io_master_0_a_bits_size;
  assign TLBuffer_4_io_in_0_a_bits_source = tile_io_master_0_a_bits_source;
  assign TLBuffer_4_io_in_0_a_bits_address = tile_io_master_0_a_bits_address;
  assign TLBuffer_4_io_in_0_a_bits_mask = tile_io_master_0_a_bits_mask;
  assign TLBuffer_4_io_in_0_a_bits_data = tile_io_master_0_a_bits_data;
  assign TLBuffer_4_io_in_0_d_ready = tile_io_master_0_d_ready;
  assign TLBuffer_4_io_out_0_a_ready = TLFIFOFixer_io_in_0_a_ready;
  assign TLBuffer_4_io_out_0_d_valid = TLFIFOFixer_io_in_0_d_valid;
  assign TLBuffer_4_io_out_0_d_bits_opcode = TLFIFOFixer_io_in_0_d_bits_opcode;
  assign TLBuffer_4_io_out_0_d_bits_size = TLFIFOFixer_io_in_0_d_bits_size;
  assign TLBuffer_4_io_out_0_d_bits_source = TLFIFOFixer_io_in_0_d_bits_source;
  assign TLBuffer_4_io_out_0_d_bits_data = TLFIFOFixer_io_in_0_d_bits_data;
  assign TLBuffer_4_io_out_0_d_bits_error = TLFIFOFixer_io_in_0_d_bits_error;
  assign IntXbar_1_io_in_0_0 = debug_1_io_debugInterrupts_0_0;
  assign IntXbar_2_io_in_1_0 = plic_io_harts_0_0;
  assign IntXbar_2_io_in_0_0 = clint_io_int_0_0;
  assign IntXbar_2_io_in_0_1 = clint_io_int_0_1;
  assign IntXing_clock = clock;
  assign IntXing_io_in_0_0 = _T_164;
  assign IntXing_io_in_0_1 = _T_165;
  assign TLToAXI4_clock = clock;
  assign TLToAXI4_reset = reset;
  assign TLToAXI4_io_in_0_a_valid = TLWidthWidget_io_out_1_a_valid;
  assign TLToAXI4_io_in_0_a_bits_opcode = TLWidthWidget_io_out_1_a_bits_opcode;
  assign TLToAXI4_io_in_0_a_bits_size = TLWidthWidget_io_out_1_a_bits_size;
  assign TLToAXI4_io_in_0_a_bits_source = TLWidthWidget_io_out_1_a_bits_source;
  assign TLToAXI4_io_in_0_a_bits_address = TLWidthWidget_io_out_1_a_bits_address;
  assign TLToAXI4_io_in_0_a_bits_mask = TLWidthWidget_io_out_1_a_bits_mask;
  assign TLToAXI4_io_in_0_a_bits_data = TLWidthWidget_io_out_1_a_bits_data;
  assign TLToAXI4_io_in_0_d_ready = TLWidthWidget_io_out_1_d_ready;
  assign TLToAXI4_io_out_0_aw_ready = AXI4IdIndexer_io_in_0_aw_ready;
  assign TLToAXI4_io_out_0_w_ready = AXI4IdIndexer_io_in_0_w_ready;
  assign TLToAXI4_io_out_0_b_valid = AXI4IdIndexer_io_in_0_b_valid;
  assign TLToAXI4_io_out_0_b_bits_id = AXI4IdIndexer_io_in_0_b_bits_id;
  assign TLToAXI4_io_out_0_b_bits_resp = AXI4IdIndexer_io_in_0_b_bits_resp;
  assign TLToAXI4_io_out_0_b_bits_user = AXI4IdIndexer_io_in_0_b_bits_user;
  assign TLToAXI4_io_out_0_ar_ready = AXI4IdIndexer_io_in_0_ar_ready;
  assign TLToAXI4_io_out_0_r_valid = AXI4IdIndexer_io_in_0_r_valid;
  assign TLToAXI4_io_out_0_r_bits_id = AXI4IdIndexer_io_in_0_r_bits_id;
  assign TLToAXI4_io_out_0_r_bits_data = AXI4IdIndexer_io_in_0_r_bits_data;
  assign TLToAXI4_io_out_0_r_bits_resp = AXI4IdIndexer_io_in_0_r_bits_resp;
  assign TLToAXI4_io_out_0_r_bits_user = AXI4IdIndexer_io_in_0_r_bits_user;
  assign TLToAXI4_io_out_0_r_bits_last = AXI4IdIndexer_io_in_0_r_bits_last;
  assign AXI4IdIndexer_io_in_0_aw_valid = TLToAXI4_io_out_0_aw_valid;
  assign AXI4IdIndexer_io_in_0_aw_bits_id = TLToAXI4_io_out_0_aw_bits_id;
  assign AXI4IdIndexer_io_in_0_aw_bits_addr = TLToAXI4_io_out_0_aw_bits_addr;
  assign AXI4IdIndexer_io_in_0_aw_bits_len = TLToAXI4_io_out_0_aw_bits_len;
  assign AXI4IdIndexer_io_in_0_aw_bits_size = TLToAXI4_io_out_0_aw_bits_size;
  assign AXI4IdIndexer_io_in_0_aw_bits_burst = TLToAXI4_io_out_0_aw_bits_burst;
  assign AXI4IdIndexer_io_in_0_aw_bits_user = TLToAXI4_io_out_0_aw_bits_user;
  assign AXI4IdIndexer_io_in_0_w_valid = TLToAXI4_io_out_0_w_valid;
  assign AXI4IdIndexer_io_in_0_w_bits_data = TLToAXI4_io_out_0_w_bits_data;
  assign AXI4IdIndexer_io_in_0_w_bits_strb = TLToAXI4_io_out_0_w_bits_strb;
  assign AXI4IdIndexer_io_in_0_w_bits_last = TLToAXI4_io_out_0_w_bits_last;
  assign AXI4IdIndexer_io_in_0_b_ready = TLToAXI4_io_out_0_b_ready;
  assign AXI4IdIndexer_io_in_0_ar_valid = TLToAXI4_io_out_0_ar_valid;
  assign AXI4IdIndexer_io_in_0_ar_bits_id = TLToAXI4_io_out_0_ar_bits_id;
  assign AXI4IdIndexer_io_in_0_ar_bits_addr = TLToAXI4_io_out_0_ar_bits_addr;
  assign AXI4IdIndexer_io_in_0_ar_bits_len = TLToAXI4_io_out_0_ar_bits_len;
  assign AXI4IdIndexer_io_in_0_ar_bits_size = TLToAXI4_io_out_0_ar_bits_size;
  assign AXI4IdIndexer_io_in_0_ar_bits_burst = TLToAXI4_io_out_0_ar_bits_burst;
  assign AXI4IdIndexer_io_in_0_ar_bits_user = TLToAXI4_io_out_0_ar_bits_user;
  assign AXI4IdIndexer_io_in_0_r_ready = TLToAXI4_io_out_0_r_ready;
  assign AXI4IdIndexer_io_out_0_aw_ready = AXI4Deinterleaver_io_in_0_aw_ready;
  assign AXI4IdIndexer_io_out_0_w_ready = AXI4Deinterleaver_io_in_0_w_ready;
  assign AXI4IdIndexer_io_out_0_b_valid = AXI4Deinterleaver_io_in_0_b_valid;
  assign AXI4IdIndexer_io_out_0_b_bits_id = AXI4Deinterleaver_io_in_0_b_bits_id;
  assign AXI4IdIndexer_io_out_0_b_bits_resp = AXI4Deinterleaver_io_in_0_b_bits_resp;
  assign AXI4IdIndexer_io_out_0_b_bits_user = AXI4Deinterleaver_io_in_0_b_bits_user;
  assign AXI4IdIndexer_io_out_0_ar_ready = AXI4Deinterleaver_io_in_0_ar_ready;
  assign AXI4IdIndexer_io_out_0_r_valid = AXI4Deinterleaver_io_in_0_r_valid;
  assign AXI4IdIndexer_io_out_0_r_bits_id = AXI4Deinterleaver_io_in_0_r_bits_id;
  assign AXI4IdIndexer_io_out_0_r_bits_data = AXI4Deinterleaver_io_in_0_r_bits_data;
  assign AXI4IdIndexer_io_out_0_r_bits_resp = AXI4Deinterleaver_io_in_0_r_bits_resp;
  assign AXI4IdIndexer_io_out_0_r_bits_user = AXI4Deinterleaver_io_in_0_r_bits_user;
  assign AXI4IdIndexer_io_out_0_r_bits_last = AXI4Deinterleaver_io_in_0_r_bits_last;
  assign AXI4Deinterleaver_clock = clock;
  assign AXI4Deinterleaver_reset = reset;
  assign AXI4Deinterleaver_io_in_0_aw_valid = AXI4IdIndexer_io_out_0_aw_valid;
  assign AXI4Deinterleaver_io_in_0_aw_bits_id = AXI4IdIndexer_io_out_0_aw_bits_id;
  assign AXI4Deinterleaver_io_in_0_aw_bits_addr = AXI4IdIndexer_io_out_0_aw_bits_addr;
  assign AXI4Deinterleaver_io_in_0_aw_bits_len = AXI4IdIndexer_io_out_0_aw_bits_len;
  assign AXI4Deinterleaver_io_in_0_aw_bits_size = AXI4IdIndexer_io_out_0_aw_bits_size;
  assign AXI4Deinterleaver_io_in_0_aw_bits_burst = AXI4IdIndexer_io_out_0_aw_bits_burst;
  assign AXI4Deinterleaver_io_in_0_aw_bits_user = AXI4IdIndexer_io_out_0_aw_bits_user;
  assign AXI4Deinterleaver_io_in_0_w_valid = AXI4IdIndexer_io_out_0_w_valid;
  assign AXI4Deinterleaver_io_in_0_w_bits_data = AXI4IdIndexer_io_out_0_w_bits_data;
  assign AXI4Deinterleaver_io_in_0_w_bits_strb = AXI4IdIndexer_io_out_0_w_bits_strb;
  assign AXI4Deinterleaver_io_in_0_w_bits_last = AXI4IdIndexer_io_out_0_w_bits_last;
  assign AXI4Deinterleaver_io_in_0_b_ready = AXI4IdIndexer_io_out_0_b_ready;
  assign AXI4Deinterleaver_io_in_0_ar_valid = AXI4IdIndexer_io_out_0_ar_valid;
  assign AXI4Deinterleaver_io_in_0_ar_bits_id = AXI4IdIndexer_io_out_0_ar_bits_id;
  assign AXI4Deinterleaver_io_in_0_ar_bits_addr = AXI4IdIndexer_io_out_0_ar_bits_addr;
  assign AXI4Deinterleaver_io_in_0_ar_bits_len = AXI4IdIndexer_io_out_0_ar_bits_len;
  assign AXI4Deinterleaver_io_in_0_ar_bits_size = AXI4IdIndexer_io_out_0_ar_bits_size;
  assign AXI4Deinterleaver_io_in_0_ar_bits_burst = AXI4IdIndexer_io_out_0_ar_bits_burst;
  assign AXI4Deinterleaver_io_in_0_ar_bits_user = AXI4IdIndexer_io_out_0_ar_bits_user;
  assign AXI4Deinterleaver_io_in_0_r_ready = AXI4IdIndexer_io_out_0_r_ready;
  assign AXI4Deinterleaver_io_out_0_aw_ready = AXI4UserYanker_io_in_0_aw_ready;
  assign AXI4Deinterleaver_io_out_0_w_ready = AXI4UserYanker_io_in_0_w_ready;
  assign AXI4Deinterleaver_io_out_0_b_valid = AXI4UserYanker_io_in_0_b_valid;
  assign AXI4Deinterleaver_io_out_0_b_bits_id = AXI4UserYanker_io_in_0_b_bits_id;
  assign AXI4Deinterleaver_io_out_0_b_bits_resp = AXI4UserYanker_io_in_0_b_bits_resp;
  assign AXI4Deinterleaver_io_out_0_b_bits_user = AXI4UserYanker_io_in_0_b_bits_user;
  assign AXI4Deinterleaver_io_out_0_ar_ready = AXI4UserYanker_io_in_0_ar_ready;
  assign AXI4Deinterleaver_io_out_0_r_valid = AXI4UserYanker_io_in_0_r_valid;
  assign AXI4Deinterleaver_io_out_0_r_bits_id = AXI4UserYanker_io_in_0_r_bits_id;
  assign AXI4Deinterleaver_io_out_0_r_bits_data = AXI4UserYanker_io_in_0_r_bits_data;
  assign AXI4Deinterleaver_io_out_0_r_bits_resp = AXI4UserYanker_io_in_0_r_bits_resp;
  assign AXI4Deinterleaver_io_out_0_r_bits_user = AXI4UserYanker_io_in_0_r_bits_user;
  assign AXI4Deinterleaver_io_out_0_r_bits_last = AXI4UserYanker_io_in_0_r_bits_last;
  assign AXI4UserYanker_clock = clock;
  assign AXI4UserYanker_reset = reset;
  assign AXI4UserYanker_io_in_0_aw_valid = AXI4Deinterleaver_io_out_0_aw_valid;
  assign AXI4UserYanker_io_in_0_aw_bits_id = AXI4Deinterleaver_io_out_0_aw_bits_id;
  assign AXI4UserYanker_io_in_0_aw_bits_addr = AXI4Deinterleaver_io_out_0_aw_bits_addr;
  assign AXI4UserYanker_io_in_0_aw_bits_len = AXI4Deinterleaver_io_out_0_aw_bits_len;
  assign AXI4UserYanker_io_in_0_aw_bits_size = AXI4Deinterleaver_io_out_0_aw_bits_size;
  assign AXI4UserYanker_io_in_0_aw_bits_burst = AXI4Deinterleaver_io_out_0_aw_bits_burst;
  assign AXI4UserYanker_io_in_0_aw_bits_user = AXI4Deinterleaver_io_out_0_aw_bits_user;
  assign AXI4UserYanker_io_in_0_w_valid = AXI4Deinterleaver_io_out_0_w_valid;
  assign AXI4UserYanker_io_in_0_w_bits_data = AXI4Deinterleaver_io_out_0_w_bits_data;
  assign AXI4UserYanker_io_in_0_w_bits_strb = AXI4Deinterleaver_io_out_0_w_bits_strb;
  assign AXI4UserYanker_io_in_0_w_bits_last = AXI4Deinterleaver_io_out_0_w_bits_last;
  assign AXI4UserYanker_io_in_0_b_ready = AXI4Deinterleaver_io_out_0_b_ready;
  assign AXI4UserYanker_io_in_0_ar_valid = AXI4Deinterleaver_io_out_0_ar_valid;
  assign AXI4UserYanker_io_in_0_ar_bits_id = AXI4Deinterleaver_io_out_0_ar_bits_id;
  assign AXI4UserYanker_io_in_0_ar_bits_addr = AXI4Deinterleaver_io_out_0_ar_bits_addr;
  assign AXI4UserYanker_io_in_0_ar_bits_len = AXI4Deinterleaver_io_out_0_ar_bits_len;
  assign AXI4UserYanker_io_in_0_ar_bits_size = AXI4Deinterleaver_io_out_0_ar_bits_size;
  assign AXI4UserYanker_io_in_0_ar_bits_burst = AXI4Deinterleaver_io_out_0_ar_bits_burst;
  assign AXI4UserYanker_io_in_0_ar_bits_user = AXI4Deinterleaver_io_out_0_ar_bits_user;
  assign AXI4UserYanker_io_in_0_r_ready = AXI4Deinterleaver_io_out_0_r_ready;
  assign AXI4UserYanker_io_out_0_aw_ready = AXI4Buffer_io_in_0_aw_ready;
  assign AXI4UserYanker_io_out_0_w_ready = AXI4Buffer_io_in_0_w_ready;
  assign AXI4UserYanker_io_out_0_b_valid = AXI4Buffer_io_in_0_b_valid;
  assign AXI4UserYanker_io_out_0_b_bits_id = AXI4Buffer_io_in_0_b_bits_id;
  assign AXI4UserYanker_io_out_0_b_bits_resp = AXI4Buffer_io_in_0_b_bits_resp;
  assign AXI4UserYanker_io_out_0_ar_ready = AXI4Buffer_io_in_0_ar_ready;
  assign AXI4UserYanker_io_out_0_r_valid = AXI4Buffer_io_in_0_r_valid;
  assign AXI4UserYanker_io_out_0_r_bits_id = AXI4Buffer_io_in_0_r_bits_id;
  assign AXI4UserYanker_io_out_0_r_bits_data = AXI4Buffer_io_in_0_r_bits_data;
  assign AXI4UserYanker_io_out_0_r_bits_resp = AXI4Buffer_io_in_0_r_bits_resp;
  assign AXI4UserYanker_io_out_0_r_bits_last = AXI4Buffer_io_in_0_r_bits_last;
  assign AXI4Buffer_clock = clock;
  assign AXI4Buffer_reset = reset;
  assign AXI4Buffer_io_in_0_aw_valid = AXI4UserYanker_io_out_0_aw_valid;
  assign AXI4Buffer_io_in_0_aw_bits_id = AXI4UserYanker_io_out_0_aw_bits_id;
  assign AXI4Buffer_io_in_0_aw_bits_addr = AXI4UserYanker_io_out_0_aw_bits_addr;
  assign AXI4Buffer_io_in_0_aw_bits_len = AXI4UserYanker_io_out_0_aw_bits_len;
  assign AXI4Buffer_io_in_0_aw_bits_size = AXI4UserYanker_io_out_0_aw_bits_size;
  assign AXI4Buffer_io_in_0_aw_bits_burst = AXI4UserYanker_io_out_0_aw_bits_burst;
  assign AXI4Buffer_io_in_0_w_valid = AXI4UserYanker_io_out_0_w_valid;
  assign AXI4Buffer_io_in_0_w_bits_data = AXI4UserYanker_io_out_0_w_bits_data;
  assign AXI4Buffer_io_in_0_w_bits_strb = AXI4UserYanker_io_out_0_w_bits_strb;
  assign AXI4Buffer_io_in_0_w_bits_last = AXI4UserYanker_io_out_0_w_bits_last;
  assign AXI4Buffer_io_in_0_b_ready = AXI4UserYanker_io_out_0_b_ready;
  assign AXI4Buffer_io_in_0_ar_valid = AXI4UserYanker_io_out_0_ar_valid;
  assign AXI4Buffer_io_in_0_ar_bits_id = AXI4UserYanker_io_out_0_ar_bits_id;
  assign AXI4Buffer_io_in_0_ar_bits_addr = AXI4UserYanker_io_out_0_ar_bits_addr;
  assign AXI4Buffer_io_in_0_ar_bits_len = AXI4UserYanker_io_out_0_ar_bits_len;
  assign AXI4Buffer_io_in_0_ar_bits_size = AXI4UserYanker_io_out_0_ar_bits_size;
  assign AXI4Buffer_io_in_0_ar_bits_burst = AXI4UserYanker_io_out_0_ar_bits_burst;
  assign AXI4Buffer_io_in_0_r_ready = AXI4UserYanker_io_out_0_r_ready;
  assign AXI4Buffer_io_out_0_aw_ready = mmio_axi4_0_aw_ready;
  assign AXI4Buffer_io_out_0_w_ready = mmio_axi4_0_w_ready;
  assign AXI4Buffer_io_out_0_b_valid = mmio_axi4_0_b_valid;
  assign AXI4Buffer_io_out_0_b_bits_id = mmio_axi4_0_b_bits_id;
  assign AXI4Buffer_io_out_0_b_bits_resp = mmio_axi4_0_b_bits_resp;
  assign AXI4Buffer_io_out_0_ar_ready = mmio_axi4_0_ar_ready;
  assign AXI4Buffer_io_out_0_r_valid = mmio_axi4_0_r_valid;
  assign AXI4Buffer_io_out_0_r_bits_id = mmio_axi4_0_r_bits_id;
  assign AXI4Buffer_io_out_0_r_bits_data = mmio_axi4_0_r_bits_data;
  assign AXI4Buffer_io_out_0_r_bits_resp = mmio_axi4_0_r_bits_resp;
  assign AXI4Buffer_io_out_0_r_bits_last = mmio_axi4_0_r_bits_last;
  assign TLBuffer_5_clock = clock;
  assign TLBuffer_5_reset = reset;
  assign TLBuffer_5_io_in_0_a_valid = TLWidthWidget_2_io_out_0_a_valid;
  assign TLBuffer_5_io_in_0_a_bits_opcode = TLWidthWidget_2_io_out_0_a_bits_opcode;
  assign TLBuffer_5_io_in_0_a_bits_param = TLWidthWidget_2_io_out_0_a_bits_param;
  assign TLBuffer_5_io_in_0_a_bits_size = TLWidthWidget_2_io_out_0_a_bits_size;
  assign TLBuffer_5_io_in_0_a_bits_source = TLWidthWidget_2_io_out_0_a_bits_source;
  assign TLBuffer_5_io_in_0_a_bits_address = TLWidthWidget_2_io_out_0_a_bits_address;
  assign TLBuffer_5_io_in_0_a_bits_mask = TLWidthWidget_2_io_out_0_a_bits_mask;
  assign TLBuffer_5_io_in_0_a_bits_data = TLWidthWidget_2_io_out_0_a_bits_data;
  assign TLBuffer_5_io_in_0_d_ready = TLWidthWidget_2_io_out_0_d_ready;
  assign TLBuffer_5_io_out_0_a_ready = TLFIFOFixer_1_io_in_0_a_ready;
  assign TLBuffer_5_io_out_0_d_valid = TLFIFOFixer_1_io_in_0_d_valid;
  assign TLBuffer_5_io_out_0_d_bits_opcode = TLFIFOFixer_1_io_in_0_d_bits_opcode;
  assign TLBuffer_5_io_out_0_d_bits_size = TLFIFOFixer_1_io_in_0_d_bits_size;
  assign TLBuffer_5_io_out_0_d_bits_source = TLFIFOFixer_1_io_in_0_d_bits_source;
  assign AXI4IdIndexer_1_io_in_0_aw_valid = l2_frontend_bus_axi4_0_aw_valid;
  assign AXI4IdIndexer_1_io_in_0_aw_bits_id = l2_frontend_bus_axi4_0_aw_bits_id;
  assign AXI4IdIndexer_1_io_in_0_aw_bits_addr = l2_frontend_bus_axi4_0_aw_bits_addr;
  assign AXI4IdIndexer_1_io_in_0_aw_bits_len = l2_frontend_bus_axi4_0_aw_bits_len;
  assign AXI4IdIndexer_1_io_in_0_aw_bits_size = l2_frontend_bus_axi4_0_aw_bits_size;
  assign AXI4IdIndexer_1_io_in_0_aw_bits_burst = l2_frontend_bus_axi4_0_aw_bits_burst;
  assign AXI4IdIndexer_1_io_in_0_w_valid = l2_frontend_bus_axi4_0_w_valid;
  assign AXI4IdIndexer_1_io_in_0_w_bits_data = l2_frontend_bus_axi4_0_w_bits_data;
  assign AXI4IdIndexer_1_io_in_0_w_bits_strb = l2_frontend_bus_axi4_0_w_bits_strb;
  assign AXI4IdIndexer_1_io_in_0_w_bits_last = l2_frontend_bus_axi4_0_w_bits_last;
  assign AXI4IdIndexer_1_io_in_0_b_ready = l2_frontend_bus_axi4_0_b_ready;
  assign AXI4IdIndexer_1_io_in_0_ar_valid = l2_frontend_bus_axi4_0_ar_valid;
  assign AXI4IdIndexer_1_io_in_0_ar_bits_id = l2_frontend_bus_axi4_0_ar_bits_id;
  assign AXI4IdIndexer_1_io_in_0_ar_bits_addr = l2_frontend_bus_axi4_0_ar_bits_addr;
  assign AXI4IdIndexer_1_io_in_0_ar_bits_len = l2_frontend_bus_axi4_0_ar_bits_len;
  assign AXI4IdIndexer_1_io_in_0_ar_bits_size = l2_frontend_bus_axi4_0_ar_bits_size;
  assign AXI4IdIndexer_1_io_in_0_ar_bits_burst = l2_frontend_bus_axi4_0_ar_bits_burst;
  assign AXI4IdIndexer_1_io_in_0_r_ready = l2_frontend_bus_axi4_0_r_ready;
  assign AXI4Fragmenter_clock = clock;
  assign AXI4Fragmenter_reset = reset;
  assign AXI4Fragmenter_io_in_0_aw_valid = AXI4IdIndexer_1_io_out_0_aw_valid;
  assign AXI4Fragmenter_io_in_0_aw_bits_id = AXI4IdIndexer_1_io_out_0_aw_bits_id;
  assign AXI4Fragmenter_io_in_0_aw_bits_addr = AXI4IdIndexer_1_io_out_0_aw_bits_addr;
  assign AXI4Fragmenter_io_in_0_aw_bits_len = AXI4IdIndexer_1_io_out_0_aw_bits_len;
  assign AXI4Fragmenter_io_in_0_aw_bits_size = AXI4IdIndexer_1_io_out_0_aw_bits_size;
  assign AXI4Fragmenter_io_in_0_aw_bits_burst = AXI4IdIndexer_1_io_out_0_aw_bits_burst;
  assign AXI4Fragmenter_io_in_0_aw_bits_user = AXI4IdIndexer_1_io_out_0_aw_bits_user;
  assign AXI4Fragmenter_io_in_0_w_valid = AXI4IdIndexer_1_io_out_0_w_valid;
  assign AXI4Fragmenter_io_in_0_w_bits_data = AXI4IdIndexer_1_io_out_0_w_bits_data;
  assign AXI4Fragmenter_io_in_0_w_bits_strb = AXI4IdIndexer_1_io_out_0_w_bits_strb;
  assign AXI4Fragmenter_io_in_0_w_bits_last = AXI4IdIndexer_1_io_out_0_w_bits_last;
  assign AXI4Fragmenter_io_in_0_b_ready = AXI4IdIndexer_1_io_out_0_b_ready;
  assign AXI4Fragmenter_io_in_0_ar_valid = AXI4IdIndexer_1_io_out_0_ar_valid;
  assign AXI4Fragmenter_io_in_0_ar_bits_id = AXI4IdIndexer_1_io_out_0_ar_bits_id;
  assign AXI4Fragmenter_io_in_0_ar_bits_addr = AXI4IdIndexer_1_io_out_0_ar_bits_addr;
  assign AXI4Fragmenter_io_in_0_ar_bits_len = AXI4IdIndexer_1_io_out_0_ar_bits_len;
  assign AXI4Fragmenter_io_in_0_ar_bits_size = AXI4IdIndexer_1_io_out_0_ar_bits_size;
  assign AXI4Fragmenter_io_in_0_ar_bits_burst = AXI4IdIndexer_1_io_out_0_ar_bits_burst;
  assign AXI4Fragmenter_io_in_0_ar_bits_user = AXI4IdIndexer_1_io_out_0_ar_bits_user;
  assign AXI4Fragmenter_io_in_0_r_ready = AXI4IdIndexer_1_io_out_0_r_ready;
  assign AXI4Fragmenter_io_out_0_aw_ready = AXI4UserYanker_1_io_in_0_aw_ready;
  assign AXI4Fragmenter_io_out_0_w_ready = AXI4UserYanker_1_io_in_0_w_ready;
  assign AXI4Fragmenter_io_out_0_b_bits_user = AXI4UserYanker_1_io_in_0_b_bits_user;
  assign AXI4Fragmenter_io_out_0_ar_ready = AXI4UserYanker_1_io_in_0_ar_ready;
  assign AXI4UserYanker_1_clock = clock;
  assign AXI4UserYanker_1_reset = reset;
  assign AXI4UserYanker_1_io_in_0_aw_valid = AXI4Fragmenter_io_out_0_aw_valid;
  assign AXI4UserYanker_1_io_in_0_aw_bits_id = AXI4Fragmenter_io_out_0_aw_bits_id;
  assign AXI4UserYanker_1_io_in_0_aw_bits_addr = AXI4Fragmenter_io_out_0_aw_bits_addr;
  assign AXI4UserYanker_1_io_in_0_aw_bits_len = AXI4Fragmenter_io_out_0_aw_bits_len;
  assign AXI4UserYanker_1_io_in_0_aw_bits_size = AXI4Fragmenter_io_out_0_aw_bits_size;
  assign AXI4UserYanker_1_io_in_0_aw_bits_user = AXI4Fragmenter_io_out_0_aw_bits_user;
  assign AXI4UserYanker_1_io_in_0_w_valid = AXI4Fragmenter_io_out_0_w_valid;
  assign AXI4UserYanker_1_io_in_0_w_bits_data = AXI4Fragmenter_io_out_0_w_bits_data;
  assign AXI4UserYanker_1_io_in_0_w_bits_strb = AXI4Fragmenter_io_out_0_w_bits_strb;
  assign AXI4UserYanker_1_io_in_0_w_bits_last = AXI4Fragmenter_io_out_0_w_bits_last;
  assign AXI4UserYanker_1_io_in_0_b_ready = AXI4Fragmenter_io_out_0_b_ready;
  assign AXI4UserYanker_1_io_in_0_ar_valid = AXI4Fragmenter_io_out_0_ar_valid;
  assign AXI4UserYanker_1_io_in_0_ar_bits_id = AXI4Fragmenter_io_out_0_ar_bits_id;
  assign AXI4UserYanker_1_io_in_0_ar_bits_addr = AXI4Fragmenter_io_out_0_ar_bits_addr;
  assign AXI4UserYanker_1_io_in_0_ar_bits_len = AXI4Fragmenter_io_out_0_ar_bits_len;
  assign AXI4UserYanker_1_io_in_0_ar_bits_size = AXI4Fragmenter_io_out_0_ar_bits_size;
  assign AXI4UserYanker_1_io_in_0_ar_bits_user = AXI4Fragmenter_io_out_0_ar_bits_user;
  assign AXI4UserYanker_1_io_in_0_r_ready = AXI4Fragmenter_io_out_0_r_ready;
  assign AXI4UserYanker_1_io_out_0_aw_ready = AXI4ToTL_io_in_0_aw_ready;
  assign AXI4UserYanker_1_io_out_0_w_ready = AXI4ToTL_io_in_0_w_ready;
  assign AXI4UserYanker_1_io_out_0_b_valid = AXI4ToTL_io_in_0_b_valid;
  assign AXI4UserYanker_1_io_out_0_b_bits_id = AXI4ToTL_io_in_0_b_bits_id;
  assign AXI4UserYanker_1_io_out_0_ar_ready = AXI4ToTL_io_in_0_ar_ready;
  assign AXI4UserYanker_1_io_out_0_r_valid = AXI4ToTL_io_in_0_r_valid;
  assign AXI4UserYanker_1_io_out_0_r_bits_id = AXI4ToTL_io_in_0_r_bits_id;
  assign AXI4UserYanker_1_io_out_0_r_bits_last = AXI4ToTL_io_in_0_r_bits_last;
  assign AXI4ToTL_clock = clock;
  assign AXI4ToTL_reset = reset;
  assign AXI4ToTL_io_in_0_aw_valid = AXI4UserYanker_1_io_out_0_aw_valid;
  assign AXI4ToTL_io_in_0_aw_bits_id = AXI4UserYanker_1_io_out_0_aw_bits_id;
  assign AXI4ToTL_io_in_0_aw_bits_addr = AXI4UserYanker_1_io_out_0_aw_bits_addr;
  assign AXI4ToTL_io_in_0_aw_bits_len = AXI4UserYanker_1_io_out_0_aw_bits_len;
  assign AXI4ToTL_io_in_0_aw_bits_size = AXI4UserYanker_1_io_out_0_aw_bits_size;
  assign AXI4ToTL_io_in_0_w_valid = AXI4UserYanker_1_io_out_0_w_valid;
  assign AXI4ToTL_io_in_0_w_bits_data = AXI4UserYanker_1_io_out_0_w_bits_data;
  assign AXI4ToTL_io_in_0_w_bits_strb = AXI4UserYanker_1_io_out_0_w_bits_strb;
  assign AXI4ToTL_io_in_0_w_bits_last = AXI4UserYanker_1_io_out_0_w_bits_last;
  assign AXI4ToTL_io_in_0_b_ready = AXI4UserYanker_1_io_out_0_b_ready;
  assign AXI4ToTL_io_in_0_ar_valid = AXI4UserYanker_1_io_out_0_ar_valid;
  assign AXI4ToTL_io_in_0_ar_bits_id = AXI4UserYanker_1_io_out_0_ar_bits_id;
  assign AXI4ToTL_io_in_0_ar_bits_addr = AXI4UserYanker_1_io_out_0_ar_bits_addr;
  assign AXI4ToTL_io_in_0_ar_bits_len = AXI4UserYanker_1_io_out_0_ar_bits_len;
  assign AXI4ToTL_io_in_0_ar_bits_size = AXI4UserYanker_1_io_out_0_ar_bits_size;
  assign AXI4ToTL_io_in_0_r_ready = AXI4UserYanker_1_io_out_0_r_ready;
  assign AXI4ToTL_io_out_0_a_ready = TLWidthWidget_2_io_in_0_a_ready;
  assign AXI4ToTL_io_out_0_d_valid = TLWidthWidget_2_io_in_0_d_valid;
  assign AXI4ToTL_io_out_0_d_bits_opcode = TLWidthWidget_2_io_in_0_d_bits_opcode;
  assign AXI4ToTL_io_out_0_d_bits_size = TLWidthWidget_2_io_in_0_d_bits_size;
  assign AXI4ToTL_io_out_0_d_bits_source = TLWidthWidget_2_io_in_0_d_bits_source;
  assign TLWidthWidget_2_clock = clock;
  assign TLWidthWidget_2_reset = reset;
  assign TLWidthWidget_2_io_in_0_a_valid = AXI4ToTL_io_out_0_a_valid;
  assign TLWidthWidget_2_io_in_0_a_bits_opcode = AXI4ToTL_io_out_0_a_bits_opcode;
  assign TLWidthWidget_2_io_in_0_a_bits_param = AXI4ToTL_io_out_0_a_bits_param;
  assign TLWidthWidget_2_io_in_0_a_bits_size = AXI4ToTL_io_out_0_a_bits_size;
  assign TLWidthWidget_2_io_in_0_a_bits_source = AXI4ToTL_io_out_0_a_bits_source;
  assign TLWidthWidget_2_io_in_0_a_bits_address = AXI4ToTL_io_out_0_a_bits_address;
  assign TLWidthWidget_2_io_in_0_a_bits_mask = AXI4ToTL_io_out_0_a_bits_mask;
  assign TLWidthWidget_2_io_in_0_a_bits_data = AXI4ToTL_io_out_0_a_bits_data;
  assign TLWidthWidget_2_io_in_0_d_ready = AXI4ToTL_io_out_0_d_ready;
  assign TLWidthWidget_2_io_out_0_a_ready = TLBuffer_5_io_in_0_a_ready;
  assign TLWidthWidget_2_io_out_0_d_valid = TLBuffer_5_io_in_0_d_valid;
  assign TLWidthWidget_2_io_out_0_d_bits_opcode = TLBuffer_5_io_in_0_d_bits_opcode;
  assign TLWidthWidget_2_io_out_0_d_bits_size = TLBuffer_5_io_in_0_d_bits_size;
  assign TLWidthWidget_2_io_out_0_d_bits_source = TLBuffer_5_io_in_0_d_bits_source;
  assign bootrom_io_in_0_a_valid = TLFragmenter_1_io_out_3_a_valid;
  assign bootrom_io_in_0_a_bits_size = TLFragmenter_1_io_out_3_a_bits_size;
  assign bootrom_io_in_0_a_bits_source = TLFragmenter_1_io_out_3_a_bits_source;
  assign bootrom_io_in_0_a_bits_address = TLFragmenter_1_io_out_3_a_bits_address;
  assign bootrom_io_in_0_d_ready = TLFragmenter_1_io_out_3_d_ready;
  assign error_clock = clock;
  assign error_reset = reset;
  assign error_io_in_0_a_valid = error_TLBuffer_io_out_0_a_valid;
  assign error_io_in_0_a_bits_opcode = error_TLBuffer_io_out_0_a_bits_opcode;
  assign error_io_in_0_a_bits_size = error_TLBuffer_io_out_0_a_bits_size;
  assign error_io_in_0_a_bits_source = error_TLBuffer_io_out_0_a_bits_source;
  assign error_io_in_0_c_valid = error_TLBuffer_io_out_0_c_valid;
  assign error_io_in_0_c_bits_param = error_TLBuffer_io_out_0_c_bits_param;
  assign error_io_in_0_c_bits_size = error_TLBuffer_io_out_0_c_bits_size;
  assign error_io_in_0_c_bits_source = error_TLBuffer_io_out_0_c_bits_source;
  assign error_io_in_0_d_ready = error_TLBuffer_io_out_0_d_ready;
  assign error_TLBuffer_clock = clock;
  assign error_TLBuffer_reset = reset;
  assign error_TLBuffer_io_in_0_a_valid = TLBuffer_1_io_out_2_a_valid;
  assign error_TLBuffer_io_in_0_a_bits_opcode = TLBuffer_1_io_out_2_a_bits_opcode;
  assign error_TLBuffer_io_in_0_a_bits_size = TLBuffer_1_io_out_2_a_bits_size;
  assign error_TLBuffer_io_in_0_a_bits_source = TLBuffer_1_io_out_2_a_bits_source;
  assign error_TLBuffer_io_in_0_d_ready = TLBuffer_1_io_out_2_d_ready;
  assign error_TLBuffer_io_out_0_a_ready = error_io_in_0_a_ready;
  assign error_TLBuffer_io_out_0_d_valid = error_io_in_0_d_valid;
  assign error_TLBuffer_io_out_0_d_bits_opcode = error_io_in_0_d_bits_opcode;
  assign error_TLBuffer_io_out_0_d_bits_param = error_io_in_0_d_bits_param;
  assign error_TLBuffer_io_out_0_d_bits_size = error_io_in_0_d_bits_size;
  assign error_TLBuffer_io_out_0_d_bits_source = error_io_in_0_d_bits_source;
  assign error_TLBuffer_io_out_0_d_bits_sink = error_io_in_0_d_bits_sink;
  assign error_TLBuffer_io_out_0_d_bits_data = error_io_in_0_d_bits_data;
  assign error_TLBuffer_io_out_0_d_bits_error = error_io_in_0_d_bits_error;
  assign _T_158 = value == 7'h63;
  assign _T_160 = value + 7'h1;
  assign _T_161 = _T_160[6:0];
  assign _GEN_0 = _T_158 ? 7'h0 : _T_161;
  assign _T_164 = interrupts[0];
  assign _T_165 = interrupts[1];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      value <= 7'h0;
    end else begin
      if (_T_158) begin
        value <= 7'h0;
      end else begin
        value <= _T_161;
      end
    end
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [3:0]  io_in_0_aw_bits_id,
  input  [11:0] io_in_0_aw_bits_addr,
  input         io_in_0_aw_bits_user,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [3:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output        io_in_0_b_bits_user,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [3:0]  io_in_0_ar_bits_id,
  input  [11:0] io_in_0_ar_bits_addr,
  input         io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [3:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output        io_in_0_r_bits_user,
  output        io_in_0_r_bits_last
);
  wire [8:0] mem_R0_addr;
  wire  mem_R0_en;
  wire  mem_R0_clk;
  wire [7:0] mem_R0_data_0;
  wire [7:0] mem_R0_data_1;
  wire [7:0] mem_R0_data_2;
  wire [7:0] mem_R0_data_3;
  wire [7:0] mem_R0_data_4;
  wire [7:0] mem_R0_data_5;
  wire [7:0] mem_R0_data_6;
  wire [7:0] mem_R0_data_7;
  wire [8:0] mem_W0_addr;
  wire  mem_W0_en;
  wire  mem_W0_clk;
  wire [7:0] mem_W0_data_0;
  wire [7:0] mem_W0_data_1;
  wire [7:0] mem_W0_data_2;
  wire [7:0] mem_W0_data_3;
  wire [7:0] mem_W0_data_4;
  wire [7:0] mem_W0_data_5;
  wire [7:0] mem_W0_data_6;
  wire [7:0] mem_W0_data_7;
  wire  mem_W0_mask_0;
  wire  mem_W0_mask_1;
  wire  mem_W0_mask_2;
  wire  mem_W0_mask_3;
  wire  mem_W0_mask_4;
  wire  mem_W0_mask_5;
  wire  mem_W0_mask_6;
  wire  mem_W0_mask_7;
  wire [8:0] _T_74;
  wire  _T_75;
  wire  _T_76;
  wire  _T_77;
  wire  _T_78;
  wire  _T_79;
  wire  _T_80;
  wire  _T_81;
  wire  _T_82;
  wire  _T_83;
  wire [1:0] _T_84;
  wire [1:0] _T_85;
  wire [3:0] _T_86;
  wire [1:0] _T_87;
  wire [1:0] _T_88;
  wire [2:0] _T_89;
  wire [4:0] _T_90;
  wire [8:0] r_addr;
  wire [8:0] _T_91;
  wire  _T_92;
  wire  _T_93;
  wire  _T_94;
  wire  _T_95;
  wire  _T_96;
  wire  _T_97;
  wire  _T_98;
  wire  _T_99;
  wire  _T_100;
  wire [1:0] _T_101;
  wire [1:0] _T_102;
  wire [3:0] _T_103;
  wire [1:0] _T_104;
  wire [1:0] _T_105;
  wire [2:0] _T_106;
  wire [4:0] _T_107;
  wire [8:0] w_addr;
  wire [12:0] _T_110;
  wire [12:0] _T_112;
  wire [12:0] _T_113;
  wire  r_sel0;
  wire [12:0] _T_117;
  wire [12:0] _T_119;
  wire [12:0] _T_120;
  wire  w_sel0;
  reg  w_full;
  reg [31:0] _RAND_0;
  reg [3:0] w_id;
  reg [31:0] _RAND_1;
  reg  w_user;
  reg [31:0] _RAND_2;
  reg  r_sel1;
  reg [31:0] _RAND_3;
  reg  w_sel1;
  reg [31:0] _RAND_4;
  wire  _T_126;
  wire  _GEN_0;
  wire  _T_128;
  wire  _GEN_1;
  wire [3:0] _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [7:0] _T_131;
  wire [7:0] _T_132;
  wire [7:0] _T_133;
  wire [7:0] _T_134;
  wire [7:0] _T_135;
  wire [7:0] _T_136;
  wire [7:0] _T_137;
  wire [7:0] _T_138;
  wire  _T_152;
  wire  _T_153;
  wire  _T_154;
  wire  _T_155;
  wire  _T_156;
  wire  _T_157;
  wire  _T_158;
  wire  _T_159;
  wire  _T_160;
  wire  _GEN_25;
  wire  _GEN_27;
  wire  _GEN_29;
  wire  _GEN_31;
  wire  _GEN_33;
  wire  _GEN_35;
  wire  _GEN_37;
  wire  _GEN_39;
  wire  _T_182;
  wire  _T_183;
  wire  _T_184;
  wire  _T_188;
  wire [1:0] _T_191;
  reg  r_full;
  reg [31:0] _RAND_5;
  reg [3:0] r_id;
  reg [31:0] _RAND_6;
  reg  r_user;
  reg [31:0] _RAND_7;
  wire  _T_196;
  wire  _GEN_40;
  wire  _T_198;
  wire  _GEN_41;
  wire [3:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  reg  _T_227;
  reg [31:0] _RAND_8;
  reg [7:0] _T_257_0;
  reg [31:0] _RAND_9;
  reg [7:0] _T_257_1;
  reg [31:0] _RAND_10;
  reg [7:0] _T_257_2;
  reg [31:0] _RAND_11;
  reg [7:0] _T_257_3;
  reg [31:0] _RAND_12;
  reg [7:0] _T_257_4;
  reg [31:0] _RAND_13;
  reg [7:0] _T_257_5;
  reg [31:0] _RAND_14;
  reg [7:0] _T_257_6;
  reg [31:0] _RAND_15;
  reg [7:0] _T_257_7;
  reg [31:0] _RAND_16;
  wire [7:0] _GEN_49;
  wire [7:0] _GEN_50;
  wire [7:0] _GEN_51;
  wire [7:0] _GEN_52;
  wire [7:0] _GEN_53;
  wire [7:0] _GEN_54;
  wire [7:0] _GEN_55;
  wire [7:0] _GEN_56;
  wire  _T_324;
  wire  _T_325;
  wire [1:0] _T_328;
  wire [15:0] _T_329;
  wire [15:0] _T_330;
  wire [31:0] _T_331;
  wire [15:0] _T_332;
  wire [15:0] _T_333;
  wire [31:0] _T_334;
  wire [63:0] _T_335;
  mem mem (
    .R0_addr(mem_R0_addr),
    .R0_en(mem_R0_en),
    .R0_clk(mem_R0_clk),
    .R0_data_0(mem_R0_data_0),
    .R0_data_1(mem_R0_data_1),
    .R0_data_2(mem_R0_data_2),
    .R0_data_3(mem_R0_data_3),
    .R0_data_4(mem_R0_data_4),
    .R0_data_5(mem_R0_data_5),
    .R0_data_6(mem_R0_data_6),
    .R0_data_7(mem_R0_data_7),
    .W0_addr(mem_W0_addr),
    .W0_en(mem_W0_en),
    .W0_clk(mem_W0_clk),
    .W0_data_0(mem_W0_data_0),
    .W0_data_1(mem_W0_data_1),
    .W0_data_2(mem_W0_data_2),
    .W0_data_3(mem_W0_data_3),
    .W0_data_4(mem_W0_data_4),
    .W0_data_5(mem_W0_data_5),
    .W0_data_6(mem_W0_data_6),
    .W0_data_7(mem_W0_data_7),
    .W0_mask_0(mem_W0_mask_0),
    .W0_mask_1(mem_W0_mask_1),
    .W0_mask_2(mem_W0_mask_2),
    .W0_mask_3(mem_W0_mask_3),
    .W0_mask_4(mem_W0_mask_4),
    .W0_mask_5(mem_W0_mask_5),
    .W0_mask_6(mem_W0_mask_6),
    .W0_mask_7(mem_W0_mask_7)
  );
  assign io_in_0_aw_ready = _T_184;
  assign io_in_0_w_ready = _T_188;
  assign io_in_0_b_valid = w_full;
  assign io_in_0_b_bits_id = w_id;
  assign io_in_0_b_bits_resp = _T_191;
  assign io_in_0_b_bits_user = w_user;
  assign io_in_0_ar_ready = _T_325;
  assign io_in_0_r_valid = r_full;
  assign io_in_0_r_bits_id = r_id;
  assign io_in_0_r_bits_data = _T_335;
  assign io_in_0_r_bits_resp = _T_328;
  assign io_in_0_r_bits_user = r_user;
  assign io_in_0_r_bits_last = 1'h1;
  assign mem_R0_addr = r_addr;
  assign mem_R0_en = _T_198;
  assign mem_R0_clk = clock;
  assign mem_W0_addr = w_addr;
  assign mem_W0_en = _T_152;
  assign mem_W0_clk = clock;
  assign mem_W0_data_0 = _T_131;
  assign mem_W0_data_1 = _T_132;
  assign mem_W0_data_2 = _T_133;
  assign mem_W0_data_3 = _T_134;
  assign mem_W0_data_4 = _T_135;
  assign mem_W0_data_5 = _T_136;
  assign mem_W0_data_6 = _T_137;
  assign mem_W0_data_7 = _T_138;
  assign mem_W0_mask_0 = _GEN_25;
  assign mem_W0_mask_1 = _GEN_27;
  assign mem_W0_mask_2 = _GEN_29;
  assign mem_W0_mask_3 = _GEN_31;
  assign mem_W0_mask_4 = _GEN_33;
  assign mem_W0_mask_5 = _GEN_35;
  assign mem_W0_mask_6 = _GEN_37;
  assign mem_W0_mask_7 = _GEN_39;
  assign _T_74 = io_in_0_ar_bits_addr[11:3];
  assign _T_75 = _T_74[0];
  assign _T_76 = _T_74[1];
  assign _T_77 = _T_74[2];
  assign _T_78 = _T_74[3];
  assign _T_79 = _T_74[4];
  assign _T_80 = _T_74[5];
  assign _T_81 = _T_74[6];
  assign _T_82 = _T_74[7];
  assign _T_83 = _T_74[8];
  assign _T_84 = {_T_76,_T_75};
  assign _T_85 = {_T_78,_T_77};
  assign _T_86 = {_T_85,_T_84};
  assign _T_87 = {_T_80,_T_79};
  assign _T_88 = {_T_83,_T_82};
  assign _T_89 = {_T_88,_T_81};
  assign _T_90 = {_T_89,_T_87};
  assign r_addr = {_T_90,_T_86};
  assign _T_91 = io_in_0_aw_bits_addr[11:3];
  assign _T_92 = _T_91[0];
  assign _T_93 = _T_91[1];
  assign _T_94 = _T_91[2];
  assign _T_95 = _T_91[3];
  assign _T_96 = _T_91[4];
  assign _T_97 = _T_91[5];
  assign _T_98 = _T_91[6];
  assign _T_99 = _T_91[7];
  assign _T_100 = _T_91[8];
  assign _T_101 = {_T_93,_T_92};
  assign _T_102 = {_T_95,_T_94};
  assign _T_103 = {_T_102,_T_101};
  assign _T_104 = {_T_97,_T_96};
  assign _T_105 = {_T_100,_T_99};
  assign _T_106 = {_T_105,_T_98};
  assign _T_107 = {_T_106,_T_104};
  assign w_addr = {_T_107,_T_103};
  assign _T_110 = {1'b0,$signed(io_in_0_ar_bits_addr)};
  assign _T_112 = $signed(_T_110) & $signed(-13'sh1000);
  assign _T_113 = $signed(_T_112);
  assign r_sel0 = $signed(_T_113) == $signed(13'sh0);
  assign _T_117 = {1'b0,$signed(io_in_0_aw_bits_addr)};
  assign _T_119 = $signed(_T_117) & $signed(-13'sh1000);
  assign _T_120 = $signed(_T_119);
  assign w_sel0 = $signed(_T_120) == $signed(13'sh0);
  assign _T_126 = io_in_0_b_ready & io_in_0_b_valid;
  assign _GEN_0 = _T_126 ? 1'h0 : w_full;
  assign _T_128 = io_in_0_aw_ready & io_in_0_aw_valid;
  assign _GEN_1 = _T_128 ? 1'h1 : _GEN_0;
  assign _GEN_2 = _T_128 ? io_in_0_aw_bits_id : w_id;
  assign _GEN_3 = _T_128 ? w_sel0 : w_sel1;
  assign _GEN_4 = _T_128 ? io_in_0_aw_bits_user : w_user;
  assign _T_131 = io_in_0_w_bits_data[7:0];
  assign _T_132 = io_in_0_w_bits_data[15:8];
  assign _T_133 = io_in_0_w_bits_data[23:16];
  assign _T_134 = io_in_0_w_bits_data[31:24];
  assign _T_135 = io_in_0_w_bits_data[39:32];
  assign _T_136 = io_in_0_w_bits_data[47:40];
  assign _T_137 = io_in_0_w_bits_data[55:48];
  assign _T_138 = io_in_0_w_bits_data[63:56];
  assign _T_152 = _T_128 & w_sel0;
  assign _T_153 = io_in_0_w_bits_strb[0];
  assign _T_154 = io_in_0_w_bits_strb[1];
  assign _T_155 = io_in_0_w_bits_strb[2];
  assign _T_156 = io_in_0_w_bits_strb[3];
  assign _T_157 = io_in_0_w_bits_strb[4];
  assign _T_158 = io_in_0_w_bits_strb[5];
  assign _T_159 = io_in_0_w_bits_strb[6];
  assign _T_160 = io_in_0_w_bits_strb[7];
  assign _GEN_25 = _T_152 ? _T_153 : 1'h0;
  assign _GEN_27 = _T_152 ? _T_154 : 1'h0;
  assign _GEN_29 = _T_152 ? _T_155 : 1'h0;
  assign _GEN_31 = _T_152 ? _T_156 : 1'h0;
  assign _GEN_33 = _T_152 ? _T_157 : 1'h0;
  assign _GEN_35 = _T_152 ? _T_158 : 1'h0;
  assign _GEN_37 = _T_152 ? _T_159 : 1'h0;
  assign _GEN_39 = _T_152 ? _T_160 : 1'h0;
  assign _T_182 = w_full == 1'h0;
  assign _T_183 = io_in_0_b_ready | _T_182;
  assign _T_184 = io_in_0_w_valid & _T_183;
  assign _T_188 = io_in_0_aw_valid & _T_183;
  assign _T_191 = w_sel1 ? 2'h0 : 2'h3;
  assign _T_196 = io_in_0_r_ready & io_in_0_r_valid;
  assign _GEN_40 = _T_196 ? 1'h0 : r_full;
  assign _T_198 = io_in_0_ar_ready & io_in_0_ar_valid;
  assign _GEN_41 = _T_198 ? 1'h1 : _GEN_40;
  assign _GEN_42 = _T_198 ? io_in_0_ar_bits_id : r_id;
  assign _GEN_43 = _T_198 ? r_sel0 : r_sel1;
  assign _GEN_44 = _T_198 ? io_in_0_ar_bits_user : r_user;
  assign _GEN_49 = _T_227 ? mem_R0_data_0 : _T_257_0;
  assign _GEN_50 = _T_227 ? mem_R0_data_1 : _T_257_1;
  assign _GEN_51 = _T_227 ? mem_R0_data_2 : _T_257_2;
  assign _GEN_52 = _T_227 ? mem_R0_data_3 : _T_257_3;
  assign _GEN_53 = _T_227 ? mem_R0_data_4 : _T_257_4;
  assign _GEN_54 = _T_227 ? mem_R0_data_5 : _T_257_5;
  assign _GEN_55 = _T_227 ? mem_R0_data_6 : _T_257_6;
  assign _GEN_56 = _T_227 ? mem_R0_data_7 : _T_257_7;
  assign _T_324 = r_full == 1'h0;
  assign _T_325 = io_in_0_r_ready | _T_324;
  assign _T_328 = r_sel1 ? 2'h0 : 2'h3;
  assign _T_329 = {_GEN_50,_GEN_49};
  assign _T_330 = {_GEN_52,_GEN_51};
  assign _T_331 = {_T_330,_T_329};
  assign _T_332 = {_GEN_54,_GEN_53};
  assign _T_333 = {_GEN_56,_GEN_55};
  assign _T_334 = {_T_333,_T_332};
  assign _T_335 = {_T_334,_T_331};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  w_full = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  w_id = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  w_user = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  r_sel1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  w_sel1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  r_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  r_id = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  r_user = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_227 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_257_0 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_257_1 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_257_2 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_257_3 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_257_4 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_257_5 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_257_6 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_257_7 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      w_full <= 1'h0;
    end else begin
      if (_T_128) begin
        w_full <= 1'h1;
      end else begin
        if (_T_126) begin
          w_full <= 1'h0;
        end
      end
    end
    if (_T_128) begin
      w_id <= io_in_0_aw_bits_id;
    end
    if (_T_128) begin
      w_user <= io_in_0_aw_bits_user;
    end
    if (_T_198) begin
      r_sel1 <= r_sel0;
    end
    if (_T_128) begin
      w_sel1 <= w_sel0;
    end
    if (reset) begin
      r_full <= 1'h0;
    end else begin
      if (_T_198) begin
        r_full <= 1'h1;
      end else begin
        if (_T_196) begin
          r_full <= 1'h0;
        end
      end
    end
    if (_T_198) begin
      r_id <= io_in_0_ar_bits_id;
    end
    if (_T_198) begin
      r_user <= io_in_0_ar_bits_user;
    end
    _T_227 <= _T_198;
    if (_T_227) begin
      _T_257_0 <= mem_R0_data_0;
    end
    if (_T_227) begin
      _T_257_1 <= mem_R0_data_1;
    end
    if (_T_227) begin
      _T_257_2 <= mem_R0_data_2;
    end
    if (_T_227) begin
      _T_257_3 <= mem_R0_data_3;
    end
    if (_T_227) begin
      _T_257_4 <= mem_R0_data_4;
    end
    if (_T_227) begin
      _T_257_5 <= mem_R0_data_5;
    end
    if (_T_227) begin
      _T_257_6 <= mem_R0_data_6;
    end
    if (_T_227) begin
      _T_257_7 <= mem_R0_data_7;
    end
  end
endmodule
module Queue_45(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [11:0] io_enq_bits_addr,
  input  [7:0]  io_enq_bits_len,
  input  [2:0]  io_enq_bits_size,
  input  [1:0]  io_enq_bits_burst,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [11:0] io_deq_bits_addr,
  output [7:0]  io_deq_bits_len,
  output [2:0]  io_deq_bits_size,
  output [1:0]  io_deq_bits_burst
);
  reg [3:0] ram_id [0:0];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_35_data;
  wire  ram_id__T_35_addr;
  wire [3:0] ram_id__T_26_data;
  wire  ram_id__T_26_addr;
  wire  ram_id__T_26_mask;
  wire  ram_id__T_26_en;
  reg [11:0] ram_addr [0:0];
  reg [31:0] _RAND_1;
  wire [11:0] ram_addr__T_35_data;
  wire  ram_addr__T_35_addr;
  wire [11:0] ram_addr__T_26_data;
  wire  ram_addr__T_26_addr;
  wire  ram_addr__T_26_mask;
  wire  ram_addr__T_26_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] _RAND_2;
  wire [7:0] ram_len__T_35_data;
  wire  ram_len__T_35_addr;
  wire [7:0] ram_len__T_26_data;
  wire  ram_len__T_26_addr;
  wire  ram_len__T_26_mask;
  wire  ram_len__T_26_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] _RAND_3;
  wire [2:0] ram_size__T_35_data;
  wire  ram_size__T_35_addr;
  wire [2:0] ram_size__T_26_data;
  wire  ram_size__T_26_addr;
  wire  ram_size__T_26_mask;
  wire  ram_size__T_26_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] _RAND_4;
  wire [1:0] ram_burst__T_35_data;
  wire  ram_burst__T_35_addr;
  wire [1:0] ram_burst__T_26_data;
  wire  ram_burst__T_26_addr;
  wire  ram_burst__T_26_mask;
  wire  ram_burst__T_26_en;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_18;
  wire  _T_21;
  wire  _T_23;
  wire  _T_29;
  wire  _GEN_12;
  wire  _T_31;
  wire  _GEN_13;
  wire  _GEN_14;
  wire [3:0] _GEN_15;
  wire [11:0] _GEN_16;
  wire [7:0] _GEN_17;
  wire [2:0] _GEN_18;
  wire [1:0] _GEN_19;
  wire  _GEN_24;
  wire  _GEN_25;
  assign io_enq_ready = _T_18;
  assign io_deq_valid = _GEN_13;
  assign io_deq_bits_id = _GEN_15;
  assign io_deq_bits_addr = _GEN_16;
  assign io_deq_bits_len = _GEN_17;
  assign io_deq_bits_size = _GEN_18;
  assign io_deq_bits_burst = _GEN_19;
  assign ram_id__T_35_addr = 1'h0;
  assign ram_id__T_35_data = ram_id[ram_id__T_35_addr];
  assign ram_id__T_26_data = io_enq_bits_id;
  assign ram_id__T_26_addr = 1'h0;
  assign ram_id__T_26_mask = _GEN_25;
  assign ram_id__T_26_en = _GEN_25;
  assign ram_addr__T_35_addr = 1'h0;
  assign ram_addr__T_35_data = ram_addr[ram_addr__T_35_addr];
  assign ram_addr__T_26_data = io_enq_bits_addr;
  assign ram_addr__T_26_addr = 1'h0;
  assign ram_addr__T_26_mask = _GEN_25;
  assign ram_addr__T_26_en = _GEN_25;
  assign ram_len__T_35_addr = 1'h0;
  assign ram_len__T_35_data = ram_len[ram_len__T_35_addr];
  assign ram_len__T_26_data = io_enq_bits_len;
  assign ram_len__T_26_addr = 1'h0;
  assign ram_len__T_26_mask = _GEN_25;
  assign ram_len__T_26_en = _GEN_25;
  assign ram_size__T_35_addr = 1'h0;
  assign ram_size__T_35_data = ram_size[ram_size__T_35_addr];
  assign ram_size__T_26_data = io_enq_bits_size;
  assign ram_size__T_26_addr = 1'h0;
  assign ram_size__T_26_mask = _GEN_25;
  assign ram_size__T_26_en = _GEN_25;
  assign ram_burst__T_35_addr = 1'h0;
  assign ram_burst__T_35_data = ram_burst[ram_burst__T_35_addr];
  assign ram_burst__T_26_data = io_enq_bits_burst;
  assign ram_burst__T_26_addr = 1'h0;
  assign ram_burst__T_26_mask = _GEN_25;
  assign ram_burst__T_26_en = _GEN_25;
  assign _T_18 = maybe_full == 1'h0;
  assign _T_21 = io_enq_ready & io_enq_valid;
  assign _T_23 = io_deq_ready & io_deq_valid;
  assign _T_29 = _GEN_25 != _GEN_24;
  assign _GEN_12 = _T_29 ? _GEN_25 : maybe_full;
  assign _T_31 = _T_18 == 1'h0;
  assign _GEN_13 = io_enq_valid ? 1'h1 : _T_31;
  assign _GEN_14 = io_deq_ready ? 1'h0 : _T_21;
  assign _GEN_15 = _T_18 ? io_enq_bits_id : ram_id__T_35_data;
  assign _GEN_16 = _T_18 ? io_enq_bits_addr : ram_addr__T_35_data;
  assign _GEN_17 = _T_18 ? io_enq_bits_len : ram_len__T_35_data;
  assign _GEN_18 = _T_18 ? io_enq_bits_size : ram_size__T_35_data;
  assign _GEN_19 = _T_18 ? io_enq_bits_burst : ram_burst__T_35_data;
  assign _GEN_24 = _T_18 ? 1'h0 : _T_23;
  assign _GEN_25 = _T_18 ? _GEN_14 : _T_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = _RAND_3[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = _RAND_4[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_26_en & ram_id__T_26_mask) begin
      ram_id[ram_id__T_26_addr] <= ram_id__T_26_data;
    end
    if(ram_addr__T_26_en & ram_addr__T_26_mask) begin
      ram_addr[ram_addr__T_26_addr] <= ram_addr__T_26_data;
    end
    if(ram_len__T_26_en & ram_len__T_26_mask) begin
      ram_len[ram_len__T_26_addr] <= ram_len__T_26_data;
    end
    if(ram_size__T_26_en & ram_size__T_26_mask) begin
      ram_size[ram_size__T_26_addr] <= ram_size__T_26_data;
    end
    if(ram_burst__T_26_en & ram_burst__T_26_mask) begin
      ram_burst[ram_burst__T_26_addr] <= ram_burst__T_26_data;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_18) begin
          if (io_deq_ready) begin
            maybe_full <= 1'h0;
          end else begin
            maybe_full <= _T_21;
          end
        end else begin
          maybe_full <= _T_21;
        end
      end
    end
  end
endmodule
module AXI4Fragmenter_1(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [3:0]  io_in_0_aw_bits_id,
  input  [11:0] io_in_0_aw_bits_addr,
  input  [7:0]  io_in_0_aw_bits_len,
  input  [2:0]  io_in_0_aw_bits_size,
  input  [1:0]  io_in_0_aw_bits_burst,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [3:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [3:0]  io_in_0_ar_bits_id,
  input  [11:0] io_in_0_ar_bits_addr,
  input  [7:0]  io_in_0_ar_bits_len,
  input  [2:0]  io_in_0_ar_bits_size,
  input  [1:0]  io_in_0_ar_bits_burst,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [3:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output        io_in_0_r_bits_last,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [3:0]  io_out_0_aw_bits_id,
  output [11:0] io_out_0_aw_bits_addr,
  output        io_out_0_aw_bits_user,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_w_bits_last,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [3:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input         io_out_0_b_bits_user,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [3:0]  io_out_0_ar_bits_id,
  output [11:0] io_out_0_ar_bits_addr,
  output        io_out_0_ar_bits_user,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [3:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input         io_out_0_r_bits_user,
  input         io_out_0_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [11:0] Queue_io_enq_bits_addr;
  wire [7:0] Queue_io_enq_bits_len;
  wire [2:0] Queue_io_enq_bits_size;
  wire [1:0] Queue_io_enq_bits_burst;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [11:0] Queue_io_deq_bits_addr;
  wire [7:0] Queue_io_deq_bits_len;
  wire [2:0] Queue_io_deq_bits_size;
  wire [1:0] Queue_io_deq_bits_burst;
  wire  _T_95_valid;
  wire [3:0] _T_95_bits_id;
  wire [11:0] _T_95_bits_addr;
  wire [7:0] _T_95_bits_len;
  wire [2:0] _T_95_bits_size;
  wire [1:0] _T_95_bits_burst;
  reg  _T_105;
  reg [31:0] _RAND_0;
  reg [11:0] _T_107;
  reg [31:0] _RAND_1;
  reg [7:0] _T_109;
  reg [31:0] _RAND_2;
  wire [7:0] _T_110;
  wire [11:0] _T_111;
  wire  _T_159;
  wire [8:0] _T_165;
  wire [8:0] _T_167;
  wire [15:0] _GEN_54;
  wire [15:0] _T_172;
  wire [15:0] _GEN_55;
  wire [16:0] _T_173;
  wire [15:0] _T_174;
  wire [15:0] _T_176;
  wire [22:0] _GEN_56;
  wire [22:0] _T_177;
  wire [14:0] _T_178;
  wire  _T_182;
  wire [15:0] _GEN_57;
  wire [15:0] _T_183;
  wire [11:0] _T_184;
  wire [14:0] _GEN_58;
  wire [14:0] _T_185;
  wire [14:0] _T_186;
  wire [15:0] _GEN_59;
  wire [15:0] _T_187;
  wire [15:0] _GEN_1;
  wire [15:0] _GEN_2;
  wire  _T_190;
  wire  _T_191;
  wire [11:0] _T_192;
  wire [9:0] _T_195;
  wire [2:0] _T_196;
  wire [2:0] _T_197;
  wire [11:0] _GEN_60;
  wire [11:0] _T_198;
  wire [11:0] _T_199;
  wire  _T_200;
  wire  _T_202;
  wire [8:0] _GEN_61;
  wire [9:0] _T_203;
  wire [9:0] _T_204;
  wire [8:0] _T_205;
  wire  _GEN_3;
  wire [15:0] _GEN_4;
  wire [8:0] _GEN_5;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [3:0] Queue_1_io_enq_bits_id;
  wire [11:0] Queue_1_io_enq_bits_addr;
  wire [7:0] Queue_1_io_enq_bits_len;
  wire [2:0] Queue_1_io_enq_bits_size;
  wire [1:0] Queue_1_io_enq_bits_burst;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [3:0] Queue_1_io_deq_bits_id;
  wire [11:0] Queue_1_io_deq_bits_addr;
  wire [7:0] Queue_1_io_deq_bits_len;
  wire [2:0] Queue_1_io_deq_bits_size;
  wire [1:0] Queue_1_io_deq_bits_burst;
  wire  _T_211_valid;
  wire [3:0] _T_211_bits_id;
  wire [11:0] _T_211_bits_addr;
  wire [7:0] _T_211_bits_len;
  wire [2:0] _T_211_bits_size;
  wire [1:0] _T_211_bits_burst;
  reg  _T_221;
  reg [31:0] _RAND_3;
  reg [11:0] _T_223;
  reg [31:0] _RAND_4;
  reg [7:0] _T_225;
  reg [31:0] _RAND_5;
  wire [7:0] _T_226;
  wire [11:0] _T_227;
  wire  _T_275;
  wire [15:0] _T_288;
  wire [15:0] _GEN_73;
  wire [16:0] _T_289;
  wire [15:0] _T_290;
  wire [15:0] _T_292;
  wire [22:0] _GEN_74;
  wire [22:0] _T_293;
  wire [14:0] _T_294;
  wire  _T_298;
  wire [15:0] _GEN_75;
  wire [15:0] _T_299;
  wire [11:0] _T_300;
  wire [14:0] _GEN_76;
  wire [14:0] _T_301;
  wire [14:0] _T_302;
  wire [15:0] _GEN_77;
  wire [15:0] _T_303;
  wire [15:0] _GEN_6;
  wire [15:0] _GEN_7;
  wire  _T_306;
  wire  _T_307;
  wire [11:0] _T_308;
  wire [9:0] _T_311;
  wire [2:0] _T_312;
  wire [2:0] _T_313;
  wire [11:0] _GEN_78;
  wire [11:0] _T_314;
  wire [11:0] _T_315;
  wire  _T_316;
  wire  _T_318;
  wire [8:0] _GEN_79;
  wire [9:0] _T_319;
  wire [9:0] _T_320;
  wire [8:0] _T_321;
  wire  _GEN_8;
  wire [15:0] _GEN_9;
  wire [8:0] _GEN_10;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [63:0] Queue_2_io_enq_bits_data;
  wire [7:0] Queue_2_io_enq_bits_strb;
  wire  Queue_2_io_enq_bits_last;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [63:0] Queue_2_io_deq_bits_data;
  wire [7:0] Queue_2_io_deq_bits_strb;
  wire  Queue_2_io_deq_bits_last;
  wire  _T_327_valid;
  wire [63:0] _T_327_bits_data;
  wire [7:0] _T_327_bits_strb;
  wire  _T_327_bits_last;
  reg  _T_333;
  reg [31:0] _RAND_6;
  wire  _T_338;
  wire  _GEN_11;
  wire  _T_340;
  wire  _GEN_12;
  wire  _T_342;
  wire  _T_343;
  wire  _T_345;
  wire  _T_347;
  wire  _T_348;
  reg [8:0] _T_351;
  reg [31:0] _RAND_7;
  wire  _T_353;
  wire [8:0] _T_355;
  wire [8:0] _T_356;
  wire  _T_358;
  wire  _T_359;
  wire [8:0] _GEN_80;
  wire [9:0] _T_360;
  wire [9:0] _T_361;
  wire [8:0] _T_362;
  wire  _T_365;
  wire  _T_367;
  wire  _T_368;
  wire  _T_369;
  wire  _T_371;
  wire  _T_373;
  wire  _T_374;
  wire  _T_375;
  wire  _T_379;
  wire  _T_381;
  wire  _T_383;
  wire  _T_384;
  wire  _T_385;
  wire  _T_386;
  wire  _T_388;
  wire  _T_390;
  wire  _T_392;
  wire  _T_394;
  wire  _T_395;
  reg [1:0] _T_469_0;
  reg [31:0] _RAND_8;
  reg [1:0] _T_469_1;
  reg [31:0] _RAND_9;
  reg [1:0] _T_469_2;
  reg [31:0] _RAND_10;
  reg [1:0] _T_469_3;
  reg [31:0] _RAND_11;
  reg [1:0] _T_469_4;
  reg [31:0] _RAND_12;
  reg [1:0] _T_469_5;
  reg [31:0] _RAND_13;
  reg [1:0] _T_469_6;
  reg [31:0] _RAND_14;
  reg [1:0] _T_469_7;
  reg [31:0] _RAND_15;
  reg [1:0] _T_469_8;
  reg [31:0] _RAND_16;
  reg [1:0] _T_469_9;
  reg [31:0] _RAND_17;
  reg [1:0] _T_469_10;
  reg [31:0] _RAND_18;
  reg [1:0] _T_469_11;
  reg [31:0] _RAND_19;
  reg [1:0] _T_469_12;
  reg [31:0] _RAND_20;
  reg [1:0] _T_469_13;
  reg [31:0] _RAND_21;
  reg [1:0] _T_469_14;
  reg [31:0] _RAND_22;
  reg [1:0] _T_469_15;
  reg [31:0] _RAND_23;
  wire [1:0] _GEN_13;
  wire [1:0] _GEN_14;
  wire [1:0] _GEN_15;
  wire [1:0] _GEN_16;
  wire [1:0] _GEN_17;
  wire [1:0] _GEN_18;
  wire [1:0] _GEN_19;
  wire [1:0] _GEN_20;
  wire [1:0] _GEN_21;
  wire [1:0] _GEN_22;
  wire [1:0] _GEN_23;
  wire [1:0] _GEN_24;
  wire [1:0] _GEN_25;
  wire [1:0] _GEN_26;
  wire [1:0] _GEN_27;
  wire [1:0] _T_525;
  wire [15:0] _T_528;
  wire  _T_530;
  wire  _T_531;
  wire  _T_532;
  wire  _T_533;
  wire  _T_534;
  wire  _T_535;
  wire  _T_536;
  wire  _T_537;
  wire  _T_538;
  wire  _T_539;
  wire  _T_540;
  wire  _T_541;
  wire  _T_542;
  wire  _T_543;
  wire  _T_544;
  wire  _T_545;
  wire  _T_546;
  wire  _T_547;
  wire [1:0] _T_549;
  wire [1:0] _T_550;
  wire [1:0] _GEN_28;
  wire  _T_552;
  wire [1:0] _T_554;
  wire [1:0] _T_555;
  wire [1:0] _GEN_29;
  wire  _T_557;
  wire [1:0] _T_559;
  wire [1:0] _T_560;
  wire [1:0] _GEN_30;
  wire  _T_562;
  wire [1:0] _T_564;
  wire [1:0] _T_565;
  wire [1:0] _GEN_31;
  wire  _T_567;
  wire [1:0] _T_569;
  wire [1:0] _T_570;
  wire [1:0] _GEN_32;
  wire  _T_572;
  wire [1:0] _T_574;
  wire [1:0] _T_575;
  wire [1:0] _GEN_33;
  wire  _T_577;
  wire [1:0] _T_579;
  wire [1:0] _T_580;
  wire [1:0] _GEN_34;
  wire  _T_582;
  wire [1:0] _T_584;
  wire [1:0] _T_585;
  wire [1:0] _GEN_35;
  wire  _T_587;
  wire [1:0] _T_589;
  wire [1:0] _T_590;
  wire [1:0] _GEN_36;
  wire  _T_592;
  wire [1:0] _T_594;
  wire [1:0] _T_595;
  wire [1:0] _GEN_37;
  wire  _T_597;
  wire [1:0] _T_599;
  wire [1:0] _T_600;
  wire [1:0] _GEN_38;
  wire  _T_602;
  wire [1:0] _T_604;
  wire [1:0] _T_605;
  wire [1:0] _GEN_39;
  wire  _T_607;
  wire [1:0] _T_609;
  wire [1:0] _T_610;
  wire [1:0] _GEN_40;
  wire  _T_612;
  wire [1:0] _T_614;
  wire [1:0] _T_615;
  wire [1:0] _GEN_41;
  wire  _T_617;
  wire [1:0] _T_619;
  wire [1:0] _T_620;
  wire [1:0] _GEN_42;
  wire  _T_622;
  wire [1:0] _T_624;
  wire [1:0] _T_625;
  wire [1:0] _GEN_43;
  Queue_45 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_len(Queue_io_enq_bits_len),
    .io_enq_bits_size(Queue_io_enq_bits_size),
    .io_enq_bits_burst(Queue_io_enq_bits_burst),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_len(Queue_io_deq_bits_len),
    .io_deq_bits_size(Queue_io_deq_bits_size),
    .io_deq_bits_burst(Queue_io_deq_bits_burst)
  );
  Queue_45 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_id(Queue_1_io_enq_bits_id),
    .io_enq_bits_addr(Queue_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_1_io_enq_bits_burst),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_id(Queue_1_io_deq_bits_id),
    .io_deq_bits_addr(Queue_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_1_io_deq_bits_burst)
  );
  Queue_11 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_data(Queue_2_io_enq_bits_data),
    .io_enq_bits_strb(Queue_2_io_enq_bits_strb),
    .io_enq_bits_last(Queue_2_io_enq_bits_last),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_data(Queue_2_io_deq_bits_data),
    .io_deq_bits_strb(Queue_2_io_deq_bits_strb),
    .io_deq_bits_last(Queue_2_io_deq_bits_last)
  );
  assign io_in_0_aw_ready = Queue_1_io_enq_ready;
  assign io_in_0_w_ready = Queue_2_io_enq_ready;
  assign io_in_0_b_valid = _T_392;
  assign io_in_0_b_bits_id = io_out_0_b_bits_id;
  assign io_in_0_b_bits_resp = _T_525;
  assign io_in_0_ar_ready = Queue_io_enq_ready;
  assign io_in_0_r_valid = io_out_0_r_valid;
  assign io_in_0_r_bits_id = io_out_0_r_bits_id;
  assign io_in_0_r_bits_data = io_out_0_r_bits_data;
  assign io_in_0_r_bits_resp = io_out_0_r_bits_resp;
  assign io_in_0_r_bits_last = _T_390;
  assign io_out_0_aw_valid = _T_343;
  assign io_out_0_aw_bits_id = _T_211_bits_id;
  assign io_out_0_aw_bits_addr = _T_315;
  assign io_out_0_aw_bits_user = _T_306;
  assign io_out_0_w_valid = _T_375;
  assign io_out_0_w_bits_data = _T_327_bits_data;
  assign io_out_0_w_bits_strb = _T_327_bits_strb;
  assign io_out_0_w_bits_last = _T_358;
  assign io_out_0_b_ready = _T_395;
  assign io_out_0_ar_valid = _T_95_valid;
  assign io_out_0_ar_bits_id = _T_95_bits_id;
  assign io_out_0_ar_bits_addr = _T_199;
  assign io_out_0_ar_bits_user = _T_190;
  assign io_out_0_r_ready = io_in_0_r_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_ar_valid;
  assign Queue_io_enq_bits_id = io_in_0_ar_bits_id;
  assign Queue_io_enq_bits_addr = io_in_0_ar_bits_addr;
  assign Queue_io_enq_bits_len = io_in_0_ar_bits_len;
  assign Queue_io_enq_bits_size = io_in_0_ar_bits_size;
  assign Queue_io_enq_bits_burst = io_in_0_ar_bits_burst;
  assign Queue_io_deq_ready = _T_191;
  assign _T_95_valid = Queue_io_deq_valid;
  assign _T_95_bits_id = Queue_io_deq_bits_id;
  assign _T_95_bits_addr = Queue_io_deq_bits_addr;
  assign _T_95_bits_len = Queue_io_deq_bits_len;
  assign _T_95_bits_size = Queue_io_deq_bits_size;
  assign _T_95_bits_burst = Queue_io_deq_bits_burst;
  assign _T_110 = _T_105 ? _T_109 : _T_95_bits_len;
  assign _T_111 = _T_105 ? _T_107 : _T_95_bits_addr;
  assign _T_159 = _T_95_bits_burst == 2'h0;
  assign _T_165 = 9'h0 << 1;
  assign _T_167 = _T_165 | 9'h1;
  assign _GEN_54 = {{7'd0}, _T_167};
  assign _T_172 = _GEN_54 << _T_95_bits_size;
  assign _GEN_55 = {{4'd0}, _T_111};
  assign _T_173 = _GEN_55 + _T_172;
  assign _T_174 = _T_173[15:0];
  assign _T_176 = {_T_95_bits_len,8'hff};
  assign _GEN_56 = {{7'd0}, _T_176};
  assign _T_177 = _GEN_56 << _T_95_bits_size;
  assign _T_178 = _T_177[22:8];
  assign _T_182 = _T_95_bits_burst == 2'h2;
  assign _GEN_57 = {{1'd0}, _T_178};
  assign _T_183 = _T_174 & _GEN_57;
  assign _T_184 = ~ _T_95_bits_addr;
  assign _GEN_58 = {{3'd0}, _T_184};
  assign _T_185 = _GEN_58 | _T_178;
  assign _T_186 = ~ _T_185;
  assign _GEN_59 = {{1'd0}, _T_186};
  assign _T_187 = _T_183 | _GEN_59;
  assign _GEN_1 = _T_182 ? _T_187 : _T_174;
  assign _GEN_2 = _T_159 ? {{4'd0}, _T_95_bits_addr} : _GEN_1;
  assign _T_190 = 8'h0 == _T_110;
  assign _T_191 = io_out_0_ar_ready & _T_190;
  assign _T_192 = ~ _T_111;
  assign _T_195 = 10'h7 << _T_95_bits_size;
  assign _T_196 = _T_195[2:0];
  assign _T_197 = ~ _T_196;
  assign _GEN_60 = {{9'd0}, _T_197};
  assign _T_198 = _T_192 | _GEN_60;
  assign _T_199 = ~ _T_198;
  assign _T_200 = io_out_0_ar_ready & _T_95_valid;
  assign _T_202 = _T_190 == 1'h0;
  assign _GEN_61 = {{1'd0}, _T_110};
  assign _T_203 = _GEN_61 - _T_167;
  assign _T_204 = $unsigned(_T_203);
  assign _T_205 = _T_204[8:0];
  assign _GEN_3 = _T_200 ? _T_202 : _T_105;
  assign _GEN_4 = _T_200 ? _GEN_2 : {{4'd0}, _T_107};
  assign _GEN_5 = _T_200 ? _T_205 : {{1'd0}, _T_109};
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_in_0_aw_valid;
  assign Queue_1_io_enq_bits_id = io_in_0_aw_bits_id;
  assign Queue_1_io_enq_bits_addr = io_in_0_aw_bits_addr;
  assign Queue_1_io_enq_bits_len = io_in_0_aw_bits_len;
  assign Queue_1_io_enq_bits_size = io_in_0_aw_bits_size;
  assign Queue_1_io_enq_bits_burst = io_in_0_aw_bits_burst;
  assign Queue_1_io_deq_ready = _T_307;
  assign _T_211_valid = Queue_1_io_deq_valid;
  assign _T_211_bits_id = Queue_1_io_deq_bits_id;
  assign _T_211_bits_addr = Queue_1_io_deq_bits_addr;
  assign _T_211_bits_len = Queue_1_io_deq_bits_len;
  assign _T_211_bits_size = Queue_1_io_deq_bits_size;
  assign _T_211_bits_burst = Queue_1_io_deq_bits_burst;
  assign _T_226 = _T_221 ? _T_225 : _T_211_bits_len;
  assign _T_227 = _T_221 ? _T_223 : _T_211_bits_addr;
  assign _T_275 = _T_211_bits_burst == 2'h0;
  assign _T_288 = _GEN_54 << _T_211_bits_size;
  assign _GEN_73 = {{4'd0}, _T_227};
  assign _T_289 = _GEN_73 + _T_288;
  assign _T_290 = _T_289[15:0];
  assign _T_292 = {_T_211_bits_len,8'hff};
  assign _GEN_74 = {{7'd0}, _T_292};
  assign _T_293 = _GEN_74 << _T_211_bits_size;
  assign _T_294 = _T_293[22:8];
  assign _T_298 = _T_211_bits_burst == 2'h2;
  assign _GEN_75 = {{1'd0}, _T_294};
  assign _T_299 = _T_290 & _GEN_75;
  assign _T_300 = ~ _T_211_bits_addr;
  assign _GEN_76 = {{3'd0}, _T_300};
  assign _T_301 = _GEN_76 | _T_294;
  assign _T_302 = ~ _T_301;
  assign _GEN_77 = {{1'd0}, _T_302};
  assign _T_303 = _T_299 | _GEN_77;
  assign _GEN_6 = _T_298 ? _T_303 : _T_290;
  assign _GEN_7 = _T_275 ? {{4'd0}, _T_211_bits_addr} : _GEN_6;
  assign _T_306 = 8'h0 == _T_226;
  assign _T_307 = _T_345 & _T_306;
  assign _T_308 = ~ _T_227;
  assign _T_311 = 10'h7 << _T_211_bits_size;
  assign _T_312 = _T_311[2:0];
  assign _T_313 = ~ _T_312;
  assign _GEN_78 = {{9'd0}, _T_313};
  assign _T_314 = _T_308 | _GEN_78;
  assign _T_315 = ~ _T_314;
  assign _T_316 = _T_345 & _T_211_valid;
  assign _T_318 = _T_306 == 1'h0;
  assign _GEN_79 = {{1'd0}, _T_226};
  assign _T_319 = _GEN_79 - _T_167;
  assign _T_320 = $unsigned(_T_319);
  assign _T_321 = _T_320[8:0];
  assign _GEN_8 = _T_316 ? _T_318 : _T_221;
  assign _GEN_9 = _T_316 ? _GEN_7 : {{4'd0}, _T_223};
  assign _GEN_10 = _T_316 ? _T_321 : {{1'd0}, _T_225};
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = io_in_0_w_valid;
  assign Queue_2_io_enq_bits_data = io_in_0_w_bits_data;
  assign Queue_2_io_enq_bits_strb = io_in_0_w_bits_strb;
  assign Queue_2_io_enq_bits_last = io_in_0_w_bits_last;
  assign Queue_2_io_deq_ready = _T_379;
  assign _T_327_valid = Queue_2_io_deq_valid;
  assign _T_327_bits_data = Queue_2_io_deq_bits_data;
  assign _T_327_bits_strb = Queue_2_io_deq_bits_strb;
  assign _T_327_bits_last = Queue_2_io_deq_bits_last;
  assign _T_338 = _T_348 & _T_353;
  assign _GEN_11 = _T_338 ? 1'h1 : _T_333;
  assign _T_340 = io_out_0_aw_ready & io_out_0_aw_valid;
  assign _GEN_12 = _T_340 ? 1'h0 : _GEN_11;
  assign _T_342 = _T_353 | _T_333;
  assign _T_343 = _T_211_valid & _T_342;
  assign _T_345 = io_out_0_aw_ready & _T_342;
  assign _T_347 = _T_333 == 1'h0;
  assign _T_348 = _T_211_valid & _T_347;
  assign _T_353 = _T_351 == 9'h0;
  assign _T_355 = _T_348 ? _T_167 : 9'h0;
  assign _T_356 = _T_353 ? _T_355 : _T_351;
  assign _T_358 = _T_356 == 9'h1;
  assign _T_359 = io_out_0_w_ready & io_out_0_w_valid;
  assign _GEN_80 = {{8'd0}, _T_359};
  assign _T_360 = _T_356 - _GEN_80;
  assign _T_361 = $unsigned(_T_360);
  assign _T_362 = _T_361[8:0];
  assign _T_365 = _T_359 == 1'h0;
  assign _T_367 = _T_356 != 9'h0;
  assign _T_368 = _T_365 | _T_367;
  assign _T_369 = _T_368 | reset;
  assign _T_371 = _T_369 == 1'h0;
  assign _T_373 = _T_353 == 1'h0;
  assign _T_374 = _T_373 | _T_348;
  assign _T_375 = _T_327_valid & _T_374;
  assign _T_379 = io_out_0_w_ready & _T_374;
  assign _T_381 = io_out_0_w_valid == 1'h0;
  assign _T_383 = _T_327_bits_last == 1'h0;
  assign _T_384 = _T_381 | _T_383;
  assign _T_385 = _T_384 | _T_358;
  assign _T_386 = _T_385 | reset;
  assign _T_388 = _T_386 == 1'h0;
  assign _T_390 = io_out_0_r_bits_last & io_out_0_r_bits_user;
  assign _T_392 = io_out_0_b_valid & io_out_0_b_bits_user;
  assign _T_394 = io_out_0_b_bits_user == 1'h0;
  assign _T_395 = io_in_0_b_ready | _T_394;
  assign _GEN_13 = 4'h1 == io_out_0_b_bits_id ? _T_469_1 : _T_469_0;
  assign _GEN_14 = 4'h2 == io_out_0_b_bits_id ? _T_469_2 : _GEN_13;
  assign _GEN_15 = 4'h3 == io_out_0_b_bits_id ? _T_469_3 : _GEN_14;
  assign _GEN_16 = 4'h4 == io_out_0_b_bits_id ? _T_469_4 : _GEN_15;
  assign _GEN_17 = 4'h5 == io_out_0_b_bits_id ? _T_469_5 : _GEN_16;
  assign _GEN_18 = 4'h6 == io_out_0_b_bits_id ? _T_469_6 : _GEN_17;
  assign _GEN_19 = 4'h7 == io_out_0_b_bits_id ? _T_469_7 : _GEN_18;
  assign _GEN_20 = 4'h8 == io_out_0_b_bits_id ? _T_469_8 : _GEN_19;
  assign _GEN_21 = 4'h9 == io_out_0_b_bits_id ? _T_469_9 : _GEN_20;
  assign _GEN_22 = 4'ha == io_out_0_b_bits_id ? _T_469_10 : _GEN_21;
  assign _GEN_23 = 4'hb == io_out_0_b_bits_id ? _T_469_11 : _GEN_22;
  assign _GEN_24 = 4'hc == io_out_0_b_bits_id ? _T_469_12 : _GEN_23;
  assign _GEN_25 = 4'hd == io_out_0_b_bits_id ? _T_469_13 : _GEN_24;
  assign _GEN_26 = 4'he == io_out_0_b_bits_id ? _T_469_14 : _GEN_25;
  assign _GEN_27 = 4'hf == io_out_0_b_bits_id ? _T_469_15 : _GEN_26;
  assign _T_525 = io_out_0_b_bits_resp | _GEN_27;
  assign _T_528 = 16'h1 << io_out_0_b_bits_id;
  assign _T_530 = _T_528[0];
  assign _T_531 = _T_528[1];
  assign _T_532 = _T_528[2];
  assign _T_533 = _T_528[3];
  assign _T_534 = _T_528[4];
  assign _T_535 = _T_528[5];
  assign _T_536 = _T_528[6];
  assign _T_537 = _T_528[7];
  assign _T_538 = _T_528[8];
  assign _T_539 = _T_528[9];
  assign _T_540 = _T_528[10];
  assign _T_541 = _T_528[11];
  assign _T_542 = _T_528[12];
  assign _T_543 = _T_528[13];
  assign _T_544 = _T_528[14];
  assign _T_545 = _T_528[15];
  assign _T_546 = io_out_0_b_ready & io_out_0_b_valid;
  assign _T_547 = _T_530 & _T_546;
  assign _T_549 = _T_469_0 | io_out_0_b_bits_resp;
  assign _T_550 = io_out_0_b_bits_user ? 2'h0 : _T_549;
  assign _GEN_28 = _T_547 ? _T_550 : _T_469_0;
  assign _T_552 = _T_531 & _T_546;
  assign _T_554 = _T_469_1 | io_out_0_b_bits_resp;
  assign _T_555 = io_out_0_b_bits_user ? 2'h0 : _T_554;
  assign _GEN_29 = _T_552 ? _T_555 : _T_469_1;
  assign _T_557 = _T_532 & _T_546;
  assign _T_559 = _T_469_2 | io_out_0_b_bits_resp;
  assign _T_560 = io_out_0_b_bits_user ? 2'h0 : _T_559;
  assign _GEN_30 = _T_557 ? _T_560 : _T_469_2;
  assign _T_562 = _T_533 & _T_546;
  assign _T_564 = _T_469_3 | io_out_0_b_bits_resp;
  assign _T_565 = io_out_0_b_bits_user ? 2'h0 : _T_564;
  assign _GEN_31 = _T_562 ? _T_565 : _T_469_3;
  assign _T_567 = _T_534 & _T_546;
  assign _T_569 = _T_469_4 | io_out_0_b_bits_resp;
  assign _T_570 = io_out_0_b_bits_user ? 2'h0 : _T_569;
  assign _GEN_32 = _T_567 ? _T_570 : _T_469_4;
  assign _T_572 = _T_535 & _T_546;
  assign _T_574 = _T_469_5 | io_out_0_b_bits_resp;
  assign _T_575 = io_out_0_b_bits_user ? 2'h0 : _T_574;
  assign _GEN_33 = _T_572 ? _T_575 : _T_469_5;
  assign _T_577 = _T_536 & _T_546;
  assign _T_579 = _T_469_6 | io_out_0_b_bits_resp;
  assign _T_580 = io_out_0_b_bits_user ? 2'h0 : _T_579;
  assign _GEN_34 = _T_577 ? _T_580 : _T_469_6;
  assign _T_582 = _T_537 & _T_546;
  assign _T_584 = _T_469_7 | io_out_0_b_bits_resp;
  assign _T_585 = io_out_0_b_bits_user ? 2'h0 : _T_584;
  assign _GEN_35 = _T_582 ? _T_585 : _T_469_7;
  assign _T_587 = _T_538 & _T_546;
  assign _T_589 = _T_469_8 | io_out_0_b_bits_resp;
  assign _T_590 = io_out_0_b_bits_user ? 2'h0 : _T_589;
  assign _GEN_36 = _T_587 ? _T_590 : _T_469_8;
  assign _T_592 = _T_539 & _T_546;
  assign _T_594 = _T_469_9 | io_out_0_b_bits_resp;
  assign _T_595 = io_out_0_b_bits_user ? 2'h0 : _T_594;
  assign _GEN_37 = _T_592 ? _T_595 : _T_469_9;
  assign _T_597 = _T_540 & _T_546;
  assign _T_599 = _T_469_10 | io_out_0_b_bits_resp;
  assign _T_600 = io_out_0_b_bits_user ? 2'h0 : _T_599;
  assign _GEN_38 = _T_597 ? _T_600 : _T_469_10;
  assign _T_602 = _T_541 & _T_546;
  assign _T_604 = _T_469_11 | io_out_0_b_bits_resp;
  assign _T_605 = io_out_0_b_bits_user ? 2'h0 : _T_604;
  assign _GEN_39 = _T_602 ? _T_605 : _T_469_11;
  assign _T_607 = _T_542 & _T_546;
  assign _T_609 = _T_469_12 | io_out_0_b_bits_resp;
  assign _T_610 = io_out_0_b_bits_user ? 2'h0 : _T_609;
  assign _GEN_40 = _T_607 ? _T_610 : _T_469_12;
  assign _T_612 = _T_543 & _T_546;
  assign _T_614 = _T_469_13 | io_out_0_b_bits_resp;
  assign _T_615 = io_out_0_b_bits_user ? 2'h0 : _T_614;
  assign _GEN_41 = _T_612 ? _T_615 : _T_469_13;
  assign _T_617 = _T_544 & _T_546;
  assign _T_619 = _T_469_14 | io_out_0_b_bits_resp;
  assign _T_620 = io_out_0_b_bits_user ? 2'h0 : _T_619;
  assign _GEN_42 = _T_617 ? _T_620 : _T_469_14;
  assign _T_622 = _T_545 & _T_546;
  assign _T_624 = _T_469_15 | io_out_0_b_bits_resp;
  assign _T_625 = io_out_0_b_bits_user ? 2'h0 : _T_624;
  assign _GEN_43 = _T_622 ? _T_625 : _T_469_15;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_105 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_107 = _RAND_1[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_109 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_221 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_223 = _RAND_4[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_225 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_333 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_351 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_469_0 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_469_1 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_469_2 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_469_3 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_469_4 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_469_5 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_469_6 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_469_7 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_469_8 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_469_9 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_469_10 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_469_11 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_469_12 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_469_13 = _RAND_21[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_469_14 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_469_15 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_105 <= 1'h0;
    end else begin
      if (_T_200) begin
        _T_105 <= _T_202;
      end
    end
    _T_107 <= _GEN_4[11:0];
    _T_109 <= _GEN_5[7:0];
    if (reset) begin
      _T_221 <= 1'h0;
    end else begin
      if (_T_316) begin
        _T_221 <= _T_318;
      end
    end
    _T_223 <= _GEN_9[11:0];
    _T_225 <= _GEN_10[7:0];
    if (reset) begin
      _T_333 <= 1'h0;
    end else begin
      if (_T_340) begin
        _T_333 <= 1'h0;
      end else begin
        if (_T_338) begin
          _T_333 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_351 <= 9'h0;
    end else begin
      _T_351 <= _T_362;
    end
    if (reset) begin
      _T_469_0 <= 2'h0;
    end else begin
      if (_T_547) begin
        if (io_out_0_b_bits_user) begin
          _T_469_0 <= 2'h0;
        end else begin
          _T_469_0 <= _T_549;
        end
      end
    end
    if (reset) begin
      _T_469_1 <= 2'h0;
    end else begin
      if (_T_552) begin
        if (io_out_0_b_bits_user) begin
          _T_469_1 <= 2'h0;
        end else begin
          _T_469_1 <= _T_554;
        end
      end
    end
    if (reset) begin
      _T_469_2 <= 2'h0;
    end else begin
      if (_T_557) begin
        if (io_out_0_b_bits_user) begin
          _T_469_2 <= 2'h0;
        end else begin
          _T_469_2 <= _T_559;
        end
      end
    end
    if (reset) begin
      _T_469_3 <= 2'h0;
    end else begin
      if (_T_562) begin
        if (io_out_0_b_bits_user) begin
          _T_469_3 <= 2'h0;
        end else begin
          _T_469_3 <= _T_564;
        end
      end
    end
    if (reset) begin
      _T_469_4 <= 2'h0;
    end else begin
      if (_T_567) begin
        if (io_out_0_b_bits_user) begin
          _T_469_4 <= 2'h0;
        end else begin
          _T_469_4 <= _T_569;
        end
      end
    end
    if (reset) begin
      _T_469_5 <= 2'h0;
    end else begin
      if (_T_572) begin
        if (io_out_0_b_bits_user) begin
          _T_469_5 <= 2'h0;
        end else begin
          _T_469_5 <= _T_574;
        end
      end
    end
    if (reset) begin
      _T_469_6 <= 2'h0;
    end else begin
      if (_T_577) begin
        if (io_out_0_b_bits_user) begin
          _T_469_6 <= 2'h0;
        end else begin
          _T_469_6 <= _T_579;
        end
      end
    end
    if (reset) begin
      _T_469_7 <= 2'h0;
    end else begin
      if (_T_582) begin
        if (io_out_0_b_bits_user) begin
          _T_469_7 <= 2'h0;
        end else begin
          _T_469_7 <= _T_584;
        end
      end
    end
    if (reset) begin
      _T_469_8 <= 2'h0;
    end else begin
      if (_T_587) begin
        if (io_out_0_b_bits_user) begin
          _T_469_8 <= 2'h0;
        end else begin
          _T_469_8 <= _T_589;
        end
      end
    end
    if (reset) begin
      _T_469_9 <= 2'h0;
    end else begin
      if (_T_592) begin
        if (io_out_0_b_bits_user) begin
          _T_469_9 <= 2'h0;
        end else begin
          _T_469_9 <= _T_594;
        end
      end
    end
    if (reset) begin
      _T_469_10 <= 2'h0;
    end else begin
      if (_T_597) begin
        if (io_out_0_b_bits_user) begin
          _T_469_10 <= 2'h0;
        end else begin
          _T_469_10 <= _T_599;
        end
      end
    end
    if (reset) begin
      _T_469_11 <= 2'h0;
    end else begin
      if (_T_602) begin
        if (io_out_0_b_bits_user) begin
          _T_469_11 <= 2'h0;
        end else begin
          _T_469_11 <= _T_604;
        end
      end
    end
    if (reset) begin
      _T_469_12 <= 2'h0;
    end else begin
      if (_T_607) begin
        if (io_out_0_b_bits_user) begin
          _T_469_12 <= 2'h0;
        end else begin
          _T_469_12 <= _T_609;
        end
      end
    end
    if (reset) begin
      _T_469_13 <= 2'h0;
    end else begin
      if (_T_612) begin
        if (io_out_0_b_bits_user) begin
          _T_469_13 <= 2'h0;
        end else begin
          _T_469_13 <= _T_614;
        end
      end
    end
    if (reset) begin
      _T_469_14 <= 2'h0;
    end else begin
      if (_T_617) begin
        if (io_out_0_b_bits_user) begin
          _T_469_14 <= 2'h0;
        end else begin
          _T_469_14 <= _T_619;
        end
      end
    end
    if (reset) begin
      _T_469_15 <= 2'h0;
    end else begin
      if (_T_622) begin
        if (io_out_0_b_bits_user) begin
          _T_469_15 <= 2'h0;
        end else begin
          _T_469_15 <= _T_624;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_371) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:172 assert (!out.w.fire() || w_todo =/= UInt(0)) // underflow impossible\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_371) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_388) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Fragmenter.scala:181 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_388) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Queue_48(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [11:0] io_enq_bits_addr,
  input         io_enq_bits_user,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [11:0] io_deq_bits_addr,
  output        io_deq_bits_user
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire  ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire  ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [11:0] ram_addr [0:1];
  reg [31:0] _RAND_1;
  wire [11:0] ram_addr__T_43_data;
  wire  ram_addr__T_43_addr;
  wire [11:0] ram_addr__T_29_data;
  wire  ram_addr__T_29_addr;
  wire  ram_addr__T_29_mask;
  wire  ram_addr__T_29_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_2;
  wire  ram_user__T_43_data;
  wire  ram_user__T_43_addr;
  wire  ram_user__T_29_data;
  wire  ram_user__T_29_addr;
  wire  ram_user__T_29_mask;
  wire  ram_user__T_29_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_13;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_14;
  wire  _T_38;
  wire  _GEN_15;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_addr = ram_addr__T_43_data;
  assign io_deq_bits_user = ram_user__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_addr__T_43_addr = value_1;
  assign ram_addr__T_43_data = ram_addr[ram_addr__T_43_addr];
  assign ram_addr__T_29_data = io_enq_bits_addr;
  assign ram_addr__T_29_addr = value;
  assign ram_addr__T_29_mask = _T_25;
  assign ram_addr__T_29_en = _T_25;
  assign ram_user__T_43_addr = value_1;
  assign ram_user__T_43_data = ram_user[ram_user__T_43_addr];
  assign ram_user__T_29_data = io_enq_bits_user;
  assign ram_user__T_29_addr = value;
  assign ram_user__T_29_mask = _T_25;
  assign ram_user__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_13 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_14 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_15 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_addr[initvar] = _RAND_1[11:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_addr__T_29_en & ram_addr__T_29_mask) begin
      ram_addr[ram_addr__T_29_addr] <= ram_addr__T_29_data;
    end
    if(ram_user__T_29_en & ram_user__T_29_mask) begin
      ram_user[ram_user__T_29_addr] <= ram_user__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_50(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [3:0] io_enq_bits_id,
  input  [1:0] io_enq_bits_resp,
  input        io_enq_bits_user,
  input        io_deq_ready,
  output       io_deq_valid,
  output [3:0] io_deq_bits_id,
  output [1:0] io_deq_bits_resp,
  output       io_deq_bits_user
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire  ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire  ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_1;
  wire [1:0] ram_resp__T_43_data;
  wire  ram_resp__T_43_addr;
  wire [1:0] ram_resp__T_29_data;
  wire  ram_resp__T_29_addr;
  wire  ram_resp__T_29_mask;
  wire  ram_resp__T_29_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_2;
  wire  ram_user__T_43_data;
  wire  ram_user__T_43_addr;
  wire  ram_user__T_29_data;
  wire  ram_user__T_29_addr;
  wire  ram_user__T_29_mask;
  wire  ram_user__T_29_en;
  reg  value;
  reg [31:0] _RAND_3;
  reg  value_1;
  reg [31:0] _RAND_4;
  reg  maybe_full;
  reg [31:0] _RAND_5;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_6;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_7;
  wire  _T_38;
  wire  _GEN_8;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_resp = ram_resp__T_43_data;
  assign io_deq_bits_user = ram_user__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_resp__T_43_addr = value_1;
  assign ram_resp__T_43_data = ram_resp[ram_resp__T_43_addr];
  assign ram_resp__T_29_data = io_enq_bits_resp;
  assign ram_resp__T_29_addr = value;
  assign ram_resp__T_29_mask = _T_25;
  assign ram_resp__T_29_en = _T_25;
  assign ram_user__T_43_addr = value_1;
  assign ram_user__T_43_data = ram_user[ram_user__T_43_addr];
  assign ram_user__T_29_data = io_enq_bits_user;
  assign ram_user__T_29_addr = value;
  assign ram_user__T_29_mask = _T_25;
  assign ram_user__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_6 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_7 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_8 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_1[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  value = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  value_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  maybe_full = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_resp__T_29_en & ram_resp__T_29_mask) begin
      ram_resp[ram_resp__T_29_addr] <= ram_resp__T_29_data;
    end
    if(ram_user__T_29_en & ram_user__T_29_mask) begin
      ram_user[ram_user__T_29_addr] <= ram_user__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module Queue_52(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [3:0]  io_enq_bits_id,
  input  [63:0] io_enq_bits_data,
  input  [1:0]  io_enq_bits_resp,
  input         io_enq_bits_user,
  input         io_enq_bits_last,
  input         io_deq_ready,
  output        io_deq_valid,
  output [3:0]  io_deq_bits_id,
  output [63:0] io_deq_bits_data,
  output [1:0]  io_deq_bits_resp,
  output        io_deq_bits_user,
  output        io_deq_bits_last
);
  reg [3:0] ram_id [0:1];
  reg [31:0] _RAND_0;
  wire [3:0] ram_id__T_43_data;
  wire  ram_id__T_43_addr;
  wire [3:0] ram_id__T_29_data;
  wire  ram_id__T_29_addr;
  wire  ram_id__T_29_mask;
  wire  ram_id__T_29_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] _RAND_1;
  wire [63:0] ram_data__T_43_data;
  wire  ram_data__T_43_addr;
  wire [63:0] ram_data__T_29_data;
  wire  ram_data__T_29_addr;
  wire  ram_data__T_29_mask;
  wire  ram_data__T_29_en;
  reg [1:0] ram_resp [0:1];
  reg [31:0] _RAND_2;
  wire [1:0] ram_resp__T_43_data;
  wire  ram_resp__T_43_addr;
  wire [1:0] ram_resp__T_29_data;
  wire  ram_resp__T_29_addr;
  wire  ram_resp__T_29_mask;
  wire  ram_resp__T_29_en;
  reg  ram_user [0:1];
  reg [31:0] _RAND_3;
  wire  ram_user__T_43_data;
  wire  ram_user__T_43_addr;
  wire  ram_user__T_29_data;
  wire  ram_user__T_29_addr;
  wire  ram_user__T_29_mask;
  wire  ram_user__T_29_en;
  reg  ram_last [0:1];
  reg [31:0] _RAND_4;
  wire  ram_last__T_43_data;
  wire  ram_last__T_43_addr;
  wire  ram_last__T_29_data;
  wire  ram_last__T_29_addr;
  wire  ram_last__T_29_mask;
  wire  ram_last__T_29_en;
  reg  value;
  reg [31:0] _RAND_5;
  reg  value_1;
  reg [31:0] _RAND_6;
  reg  maybe_full;
  reg [31:0] _RAND_7;
  wire  _T_20;
  wire  _T_22;
  wire  _T_23;
  wire  _T_24;
  wire  _T_25;
  wire  _T_27;
  wire [1:0] _T_32;
  wire  _T_33;
  wire  _GEN_8;
  wire [1:0] _T_36;
  wire  _T_37;
  wire  _GEN_9;
  wire  _T_38;
  wire  _GEN_10;
  wire  _T_40;
  wire  _T_42;
  assign io_enq_ready = _T_42;
  assign io_deq_valid = _T_40;
  assign io_deq_bits_id = ram_id__T_43_data;
  assign io_deq_bits_data = ram_data__T_43_data;
  assign io_deq_bits_resp = ram_resp__T_43_data;
  assign io_deq_bits_user = ram_user__T_43_data;
  assign io_deq_bits_last = ram_last__T_43_data;
  assign ram_id__T_43_addr = value_1;
  assign ram_id__T_43_data = ram_id[ram_id__T_43_addr];
  assign ram_id__T_29_data = io_enq_bits_id;
  assign ram_id__T_29_addr = value;
  assign ram_id__T_29_mask = _T_25;
  assign ram_id__T_29_en = _T_25;
  assign ram_data__T_43_addr = value_1;
  assign ram_data__T_43_data = ram_data[ram_data__T_43_addr];
  assign ram_data__T_29_data = io_enq_bits_data;
  assign ram_data__T_29_addr = value;
  assign ram_data__T_29_mask = _T_25;
  assign ram_data__T_29_en = _T_25;
  assign ram_resp__T_43_addr = value_1;
  assign ram_resp__T_43_data = ram_resp[ram_resp__T_43_addr];
  assign ram_resp__T_29_data = io_enq_bits_resp;
  assign ram_resp__T_29_addr = value;
  assign ram_resp__T_29_mask = _T_25;
  assign ram_resp__T_29_en = _T_25;
  assign ram_user__T_43_addr = value_1;
  assign ram_user__T_43_data = ram_user[ram_user__T_43_addr];
  assign ram_user__T_29_data = io_enq_bits_user;
  assign ram_user__T_29_addr = value;
  assign ram_user__T_29_mask = _T_25;
  assign ram_user__T_29_en = _T_25;
  assign ram_last__T_43_addr = value_1;
  assign ram_last__T_43_data = ram_last[ram_last__T_43_addr];
  assign ram_last__T_29_data = io_enq_bits_last;
  assign ram_last__T_29_addr = value;
  assign ram_last__T_29_mask = _T_25;
  assign ram_last__T_29_en = _T_25;
  assign _T_20 = value == value_1;
  assign _T_22 = maybe_full == 1'h0;
  assign _T_23 = _T_20 & _T_22;
  assign _T_24 = _T_20 & maybe_full;
  assign _T_25 = io_enq_ready & io_enq_valid;
  assign _T_27 = io_deq_ready & io_deq_valid;
  assign _T_32 = value + 1'h1;
  assign _T_33 = _T_32[0:0];
  assign _GEN_8 = _T_25 ? _T_33 : value;
  assign _T_36 = value_1 + 1'h1;
  assign _T_37 = _T_36[0:0];
  assign _GEN_9 = _T_27 ? _T_37 : value_1;
  assign _T_38 = _T_25 != _T_27;
  assign _GEN_10 = _T_38 ? _T_25 : maybe_full;
  assign _T_40 = _T_23 == 1'h0;
  assign _T_42 = _T_24 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = _RAND_0[3:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = _RAND_1[63:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = _RAND_2[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  value = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  value_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  maybe_full = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(ram_id__T_29_en & ram_id__T_29_mask) begin
      ram_id[ram_id__T_29_addr] <= ram_id__T_29_data;
    end
    if(ram_data__T_29_en & ram_data__T_29_mask) begin
      ram_data[ram_data__T_29_addr] <= ram_data__T_29_data;
    end
    if(ram_resp__T_29_en & ram_resp__T_29_mask) begin
      ram_resp[ram_resp__T_29_addr] <= ram_resp__T_29_data;
    end
    if(ram_user__T_29_en & ram_user__T_29_mask) begin
      ram_user[ram_user__T_29_addr] <= ram_user__T_29_data;
    end
    if(ram_last__T_29_en & ram_last__T_29_mask) begin
      ram_last[ram_last__T_29_addr] <= ram_last__T_29_data;
    end
    if (reset) begin
      value <= 1'h0;
    end else begin
      if (_T_25) begin
        value <= _T_33;
      end
    end
    if (reset) begin
      value_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        value_1 <= _T_37;
      end
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else begin
      if (_T_38) begin
        maybe_full <= _T_25;
      end
    end
  end
endmodule
module AXI4Buffer_1(
  input         clock,
  input         reset,
  output        io_in_0_aw_ready,
  input         io_in_0_aw_valid,
  input  [3:0]  io_in_0_aw_bits_id,
  input  [11:0] io_in_0_aw_bits_addr,
  input         io_in_0_aw_bits_user,
  output        io_in_0_w_ready,
  input         io_in_0_w_valid,
  input  [63:0] io_in_0_w_bits_data,
  input  [7:0]  io_in_0_w_bits_strb,
  input         io_in_0_w_bits_last,
  input         io_in_0_b_ready,
  output        io_in_0_b_valid,
  output [3:0]  io_in_0_b_bits_id,
  output [1:0]  io_in_0_b_bits_resp,
  output        io_in_0_b_bits_user,
  output        io_in_0_ar_ready,
  input         io_in_0_ar_valid,
  input  [3:0]  io_in_0_ar_bits_id,
  input  [11:0] io_in_0_ar_bits_addr,
  input         io_in_0_ar_bits_user,
  input         io_in_0_r_ready,
  output        io_in_0_r_valid,
  output [3:0]  io_in_0_r_bits_id,
  output [63:0] io_in_0_r_bits_data,
  output [1:0]  io_in_0_r_bits_resp,
  output        io_in_0_r_bits_user,
  output        io_in_0_r_bits_last,
  input         io_out_0_aw_ready,
  output        io_out_0_aw_valid,
  output [3:0]  io_out_0_aw_bits_id,
  output [11:0] io_out_0_aw_bits_addr,
  output        io_out_0_aw_bits_user,
  input         io_out_0_w_ready,
  output        io_out_0_w_valid,
  output [63:0] io_out_0_w_bits_data,
  output [7:0]  io_out_0_w_bits_strb,
  output        io_out_0_b_ready,
  input         io_out_0_b_valid,
  input  [3:0]  io_out_0_b_bits_id,
  input  [1:0]  io_out_0_b_bits_resp,
  input         io_out_0_b_bits_user,
  input         io_out_0_ar_ready,
  output        io_out_0_ar_valid,
  output [3:0]  io_out_0_ar_bits_id,
  output [11:0] io_out_0_ar_bits_addr,
  output        io_out_0_ar_bits_user,
  output        io_out_0_r_ready,
  input         io_out_0_r_valid,
  input  [3:0]  io_out_0_r_bits_id,
  input  [63:0] io_out_0_r_bits_data,
  input  [1:0]  io_out_0_r_bits_resp,
  input         io_out_0_r_bits_user,
  input         io_out_0_r_bits_last
);
  wire  Queue_clock;
  wire  Queue_reset;
  wire  Queue_io_enq_ready;
  wire  Queue_io_enq_valid;
  wire [3:0] Queue_io_enq_bits_id;
  wire [11:0] Queue_io_enq_bits_addr;
  wire  Queue_io_enq_bits_user;
  wire  Queue_io_deq_ready;
  wire  Queue_io_deq_valid;
  wire [3:0] Queue_io_deq_bits_id;
  wire [11:0] Queue_io_deq_bits_addr;
  wire  Queue_io_deq_bits_user;
  wire  _T_95_valid;
  wire [3:0] _T_95_bits_id;
  wire [11:0] _T_95_bits_addr;
  wire  _T_95_bits_user;
  wire  Queue_1_clock;
  wire  Queue_1_reset;
  wire  Queue_1_io_enq_ready;
  wire  Queue_1_io_enq_valid;
  wire [63:0] Queue_1_io_enq_bits_data;
  wire [7:0] Queue_1_io_enq_bits_strb;
  wire  Queue_1_io_enq_bits_last;
  wire  Queue_1_io_deq_ready;
  wire  Queue_1_io_deq_valid;
  wire [63:0] Queue_1_io_deq_bits_data;
  wire [7:0] Queue_1_io_deq_bits_strb;
  wire  Queue_1_io_deq_bits_last;
  wire  _T_104_valid;
  wire [63:0] _T_104_bits_data;
  wire [7:0] _T_104_bits_strb;
  wire  Queue_2_clock;
  wire  Queue_2_reset;
  wire  Queue_2_io_enq_ready;
  wire  Queue_2_io_enq_valid;
  wire [3:0] Queue_2_io_enq_bits_id;
  wire [1:0] Queue_2_io_enq_bits_resp;
  wire  Queue_2_io_enq_bits_user;
  wire  Queue_2_io_deq_ready;
  wire  Queue_2_io_deq_valid;
  wire [3:0] Queue_2_io_deq_bits_id;
  wire [1:0] Queue_2_io_deq_bits_resp;
  wire  Queue_2_io_deq_bits_user;
  wire  _T_113_valid;
  wire [3:0] _T_113_bits_id;
  wire [1:0] _T_113_bits_resp;
  wire  _T_113_bits_user;
  wire  Queue_3_clock;
  wire  Queue_3_reset;
  wire  Queue_3_io_enq_ready;
  wire  Queue_3_io_enq_valid;
  wire [3:0] Queue_3_io_enq_bits_id;
  wire [11:0] Queue_3_io_enq_bits_addr;
  wire  Queue_3_io_enq_bits_user;
  wire  Queue_3_io_deq_ready;
  wire  Queue_3_io_deq_valid;
  wire [3:0] Queue_3_io_deq_bits_id;
  wire [11:0] Queue_3_io_deq_bits_addr;
  wire  Queue_3_io_deq_bits_user;
  wire  _T_122_valid;
  wire [3:0] _T_122_bits_id;
  wire [11:0] _T_122_bits_addr;
  wire  _T_122_bits_user;
  wire  Queue_4_clock;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [3:0] Queue_4_io_enq_bits_id;
  wire [63:0] Queue_4_io_enq_bits_data;
  wire [1:0] Queue_4_io_enq_bits_resp;
  wire  Queue_4_io_enq_bits_user;
  wire  Queue_4_io_enq_bits_last;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [3:0] Queue_4_io_deq_bits_id;
  wire [63:0] Queue_4_io_deq_bits_data;
  wire [1:0] Queue_4_io_deq_bits_resp;
  wire  Queue_4_io_deq_bits_user;
  wire  Queue_4_io_deq_bits_last;
  wire  _T_131_valid;
  wire [3:0] _T_131_bits_id;
  wire [63:0] _T_131_bits_data;
  wire [1:0] _T_131_bits_resp;
  wire  _T_131_bits_user;
  wire  _T_131_bits_last;
  Queue_48 Queue (
    .clock(Queue_clock),
    .reset(Queue_reset),
    .io_enq_ready(Queue_io_enq_ready),
    .io_enq_valid(Queue_io_enq_valid),
    .io_enq_bits_id(Queue_io_enq_bits_id),
    .io_enq_bits_addr(Queue_io_enq_bits_addr),
    .io_enq_bits_user(Queue_io_enq_bits_user),
    .io_deq_ready(Queue_io_deq_ready),
    .io_deq_valid(Queue_io_deq_valid),
    .io_deq_bits_id(Queue_io_deq_bits_id),
    .io_deq_bits_addr(Queue_io_deq_bits_addr),
    .io_deq_bits_user(Queue_io_deq_bits_user)
  );
  Queue_26 Queue_1 (
    .clock(Queue_1_clock),
    .reset(Queue_1_reset),
    .io_enq_ready(Queue_1_io_enq_ready),
    .io_enq_valid(Queue_1_io_enq_valid),
    .io_enq_bits_data(Queue_1_io_enq_bits_data),
    .io_enq_bits_strb(Queue_1_io_enq_bits_strb),
    .io_enq_bits_last(Queue_1_io_enq_bits_last),
    .io_deq_ready(Queue_1_io_deq_ready),
    .io_deq_valid(Queue_1_io_deq_valid),
    .io_deq_bits_data(Queue_1_io_deq_bits_data),
    .io_deq_bits_strb(Queue_1_io_deq_bits_strb),
    .io_deq_bits_last(Queue_1_io_deq_bits_last)
  );
  Queue_50 Queue_2 (
    .clock(Queue_2_clock),
    .reset(Queue_2_reset),
    .io_enq_ready(Queue_2_io_enq_ready),
    .io_enq_valid(Queue_2_io_enq_valid),
    .io_enq_bits_id(Queue_2_io_enq_bits_id),
    .io_enq_bits_resp(Queue_2_io_enq_bits_resp),
    .io_enq_bits_user(Queue_2_io_enq_bits_user),
    .io_deq_ready(Queue_2_io_deq_ready),
    .io_deq_valid(Queue_2_io_deq_valid),
    .io_deq_bits_id(Queue_2_io_deq_bits_id),
    .io_deq_bits_resp(Queue_2_io_deq_bits_resp),
    .io_deq_bits_user(Queue_2_io_deq_bits_user)
  );
  Queue_48 Queue_3 (
    .clock(Queue_3_clock),
    .reset(Queue_3_reset),
    .io_enq_ready(Queue_3_io_enq_ready),
    .io_enq_valid(Queue_3_io_enq_valid),
    .io_enq_bits_id(Queue_3_io_enq_bits_id),
    .io_enq_bits_addr(Queue_3_io_enq_bits_addr),
    .io_enq_bits_user(Queue_3_io_enq_bits_user),
    .io_deq_ready(Queue_3_io_deq_ready),
    .io_deq_valid(Queue_3_io_deq_valid),
    .io_deq_bits_id(Queue_3_io_deq_bits_id),
    .io_deq_bits_addr(Queue_3_io_deq_bits_addr),
    .io_deq_bits_user(Queue_3_io_deq_bits_user)
  );
  Queue_52 Queue_4 (
    .clock(Queue_4_clock),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_id(Queue_4_io_enq_bits_id),
    .io_enq_bits_data(Queue_4_io_enq_bits_data),
    .io_enq_bits_resp(Queue_4_io_enq_bits_resp),
    .io_enq_bits_user(Queue_4_io_enq_bits_user),
    .io_enq_bits_last(Queue_4_io_enq_bits_last),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_id(Queue_4_io_deq_bits_id),
    .io_deq_bits_data(Queue_4_io_deq_bits_data),
    .io_deq_bits_resp(Queue_4_io_deq_bits_resp),
    .io_deq_bits_user(Queue_4_io_deq_bits_user),
    .io_deq_bits_last(Queue_4_io_deq_bits_last)
  );
  assign io_in_0_aw_ready = Queue_io_enq_ready;
  assign io_in_0_w_ready = Queue_1_io_enq_ready;
  assign io_in_0_b_valid = _T_113_valid;
  assign io_in_0_b_bits_id = _T_113_bits_id;
  assign io_in_0_b_bits_resp = _T_113_bits_resp;
  assign io_in_0_b_bits_user = _T_113_bits_user;
  assign io_in_0_ar_ready = Queue_3_io_enq_ready;
  assign io_in_0_r_valid = _T_131_valid;
  assign io_in_0_r_bits_id = _T_131_bits_id;
  assign io_in_0_r_bits_data = _T_131_bits_data;
  assign io_in_0_r_bits_resp = _T_131_bits_resp;
  assign io_in_0_r_bits_user = _T_131_bits_user;
  assign io_in_0_r_bits_last = _T_131_bits_last;
  assign io_out_0_aw_valid = _T_95_valid;
  assign io_out_0_aw_bits_id = _T_95_bits_id;
  assign io_out_0_aw_bits_addr = _T_95_bits_addr;
  assign io_out_0_aw_bits_user = _T_95_bits_user;
  assign io_out_0_w_valid = _T_104_valid;
  assign io_out_0_w_bits_data = _T_104_bits_data;
  assign io_out_0_w_bits_strb = _T_104_bits_strb;
  assign io_out_0_b_ready = Queue_2_io_enq_ready;
  assign io_out_0_ar_valid = _T_122_valid;
  assign io_out_0_ar_bits_id = _T_122_bits_id;
  assign io_out_0_ar_bits_addr = _T_122_bits_addr;
  assign io_out_0_ar_bits_user = _T_122_bits_user;
  assign io_out_0_r_ready = Queue_4_io_enq_ready;
  assign Queue_clock = clock;
  assign Queue_reset = reset;
  assign Queue_io_enq_valid = io_in_0_aw_valid;
  assign Queue_io_enq_bits_id = io_in_0_aw_bits_id;
  assign Queue_io_enq_bits_addr = io_in_0_aw_bits_addr;
  assign Queue_io_enq_bits_user = io_in_0_aw_bits_user;
  assign Queue_io_deq_ready = io_out_0_aw_ready;
  assign _T_95_valid = Queue_io_deq_valid;
  assign _T_95_bits_id = Queue_io_deq_bits_id;
  assign _T_95_bits_addr = Queue_io_deq_bits_addr;
  assign _T_95_bits_user = Queue_io_deq_bits_user;
  assign Queue_1_clock = clock;
  assign Queue_1_reset = reset;
  assign Queue_1_io_enq_valid = io_in_0_w_valid;
  assign Queue_1_io_enq_bits_data = io_in_0_w_bits_data;
  assign Queue_1_io_enq_bits_strb = io_in_0_w_bits_strb;
  assign Queue_1_io_enq_bits_last = io_in_0_w_bits_last;
  assign Queue_1_io_deq_ready = io_out_0_w_ready;
  assign _T_104_valid = Queue_1_io_deq_valid;
  assign _T_104_bits_data = Queue_1_io_deq_bits_data;
  assign _T_104_bits_strb = Queue_1_io_deq_bits_strb;
  assign Queue_2_clock = clock;
  assign Queue_2_reset = reset;
  assign Queue_2_io_enq_valid = io_out_0_b_valid;
  assign Queue_2_io_enq_bits_id = io_out_0_b_bits_id;
  assign Queue_2_io_enq_bits_resp = io_out_0_b_bits_resp;
  assign Queue_2_io_enq_bits_user = io_out_0_b_bits_user;
  assign Queue_2_io_deq_ready = io_in_0_b_ready;
  assign _T_113_valid = Queue_2_io_deq_valid;
  assign _T_113_bits_id = Queue_2_io_deq_bits_id;
  assign _T_113_bits_resp = Queue_2_io_deq_bits_resp;
  assign _T_113_bits_user = Queue_2_io_deq_bits_user;
  assign Queue_3_clock = clock;
  assign Queue_3_reset = reset;
  assign Queue_3_io_enq_valid = io_in_0_ar_valid;
  assign Queue_3_io_enq_bits_id = io_in_0_ar_bits_id;
  assign Queue_3_io_enq_bits_addr = io_in_0_ar_bits_addr;
  assign Queue_3_io_enq_bits_user = io_in_0_ar_bits_user;
  assign Queue_3_io_deq_ready = io_out_0_ar_ready;
  assign _T_122_valid = Queue_3_io_deq_valid;
  assign _T_122_bits_id = Queue_3_io_deq_bits_id;
  assign _T_122_bits_addr = Queue_3_io_deq_bits_addr;
  assign _T_122_bits_user = Queue_3_io_deq_bits_user;
  assign Queue_4_clock = clock;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = io_out_0_r_valid;
  assign Queue_4_io_enq_bits_id = io_out_0_r_bits_id;
  assign Queue_4_io_enq_bits_data = io_out_0_r_bits_data;
  assign Queue_4_io_enq_bits_resp = io_out_0_r_bits_resp;
  assign Queue_4_io_enq_bits_user = io_out_0_r_bits_user;
  assign Queue_4_io_enq_bits_last = io_out_0_r_bits_last;
  assign Queue_4_io_deq_ready = io_in_0_r_ready;
  assign _T_131_valid = Queue_4_io_deq_valid;
  assign _T_131_bits_id = Queue_4_io_deq_bits_id;
  assign _T_131_bits_data = Queue_4_io_deq_bits_data;
  assign _T_131_bits_resp = Queue_4_io_deq_bits_resp;
  assign _T_131_bits_user = Queue_4_io_deq_bits_user;
  assign _T_131_bits_last = Queue_4_io_deq_bits_last;
endmodule
module SimAXIMem(
  input         clock,
  input         reset,
  output        io_axi4_0_aw_ready,
  input         io_axi4_0_aw_valid,
  input  [3:0]  io_axi4_0_aw_bits_id,
  input  [11:0] io_axi4_0_aw_bits_addr,
  input  [7:0]  io_axi4_0_aw_bits_len,
  input  [2:0]  io_axi4_0_aw_bits_size,
  input  [1:0]  io_axi4_0_aw_bits_burst,
  output        io_axi4_0_w_ready,
  input         io_axi4_0_w_valid,
  input  [63:0] io_axi4_0_w_bits_data,
  input  [7:0]  io_axi4_0_w_bits_strb,
  input         io_axi4_0_w_bits_last,
  input         io_axi4_0_b_ready,
  output        io_axi4_0_b_valid,
  output [3:0]  io_axi4_0_b_bits_id,
  output [1:0]  io_axi4_0_b_bits_resp,
  output        io_axi4_0_ar_ready,
  input         io_axi4_0_ar_valid,
  input  [3:0]  io_axi4_0_ar_bits_id,
  input  [11:0] io_axi4_0_ar_bits_addr,
  input  [7:0]  io_axi4_0_ar_bits_len,
  input  [2:0]  io_axi4_0_ar_bits_size,
  input  [1:0]  io_axi4_0_ar_bits_burst,
  input         io_axi4_0_r_ready,
  output        io_axi4_0_r_valid,
  output [3:0]  io_axi4_0_r_bits_id,
  output [63:0] io_axi4_0_r_bits_data,
  output [1:0]  io_axi4_0_r_bits_resp,
  output        io_axi4_0_r_bits_last
);
  wire  AXI4RAM_clock;
  wire  AXI4RAM_reset;
  wire  AXI4RAM_io_in_0_aw_ready;
  wire  AXI4RAM_io_in_0_aw_valid;
  wire [3:0] AXI4RAM_io_in_0_aw_bits_id;
  wire [11:0] AXI4RAM_io_in_0_aw_bits_addr;
  wire  AXI4RAM_io_in_0_aw_bits_user;
  wire  AXI4RAM_io_in_0_w_ready;
  wire  AXI4RAM_io_in_0_w_valid;
  wire [63:0] AXI4RAM_io_in_0_w_bits_data;
  wire [7:0] AXI4RAM_io_in_0_w_bits_strb;
  wire  AXI4RAM_io_in_0_b_ready;
  wire  AXI4RAM_io_in_0_b_valid;
  wire [3:0] AXI4RAM_io_in_0_b_bits_id;
  wire [1:0] AXI4RAM_io_in_0_b_bits_resp;
  wire  AXI4RAM_io_in_0_b_bits_user;
  wire  AXI4RAM_io_in_0_ar_ready;
  wire  AXI4RAM_io_in_0_ar_valid;
  wire [3:0] AXI4RAM_io_in_0_ar_bits_id;
  wire [11:0] AXI4RAM_io_in_0_ar_bits_addr;
  wire  AXI4RAM_io_in_0_ar_bits_user;
  wire  AXI4RAM_io_in_0_r_ready;
  wire  AXI4RAM_io_in_0_r_valid;
  wire [3:0] AXI4RAM_io_in_0_r_bits_id;
  wire [63:0] AXI4RAM_io_in_0_r_bits_data;
  wire [1:0] AXI4RAM_io_in_0_r_bits_resp;
  wire  AXI4RAM_io_in_0_r_bits_user;
  wire  AXI4RAM_io_in_0_r_bits_last;
  wire  AXI4Fragmenter_clock;
  wire  AXI4Fragmenter_reset;
  wire  AXI4Fragmenter_io_in_0_aw_ready;
  wire  AXI4Fragmenter_io_in_0_aw_valid;
  wire [3:0] AXI4Fragmenter_io_in_0_aw_bits_id;
  wire [11:0] AXI4Fragmenter_io_in_0_aw_bits_addr;
  wire [7:0] AXI4Fragmenter_io_in_0_aw_bits_len;
  wire [2:0] AXI4Fragmenter_io_in_0_aw_bits_size;
  wire [1:0] AXI4Fragmenter_io_in_0_aw_bits_burst;
  wire  AXI4Fragmenter_io_in_0_w_ready;
  wire  AXI4Fragmenter_io_in_0_w_valid;
  wire [63:0] AXI4Fragmenter_io_in_0_w_bits_data;
  wire [7:0] AXI4Fragmenter_io_in_0_w_bits_strb;
  wire  AXI4Fragmenter_io_in_0_w_bits_last;
  wire  AXI4Fragmenter_io_in_0_b_ready;
  wire  AXI4Fragmenter_io_in_0_b_valid;
  wire [3:0] AXI4Fragmenter_io_in_0_b_bits_id;
  wire [1:0] AXI4Fragmenter_io_in_0_b_bits_resp;
  wire  AXI4Fragmenter_io_in_0_ar_ready;
  wire  AXI4Fragmenter_io_in_0_ar_valid;
  wire [3:0] AXI4Fragmenter_io_in_0_ar_bits_id;
  wire [11:0] AXI4Fragmenter_io_in_0_ar_bits_addr;
  wire [7:0] AXI4Fragmenter_io_in_0_ar_bits_len;
  wire [2:0] AXI4Fragmenter_io_in_0_ar_bits_size;
  wire [1:0] AXI4Fragmenter_io_in_0_ar_bits_burst;
  wire  AXI4Fragmenter_io_in_0_r_ready;
  wire  AXI4Fragmenter_io_in_0_r_valid;
  wire [3:0] AXI4Fragmenter_io_in_0_r_bits_id;
  wire [63:0] AXI4Fragmenter_io_in_0_r_bits_data;
  wire [1:0] AXI4Fragmenter_io_in_0_r_bits_resp;
  wire  AXI4Fragmenter_io_in_0_r_bits_last;
  wire  AXI4Fragmenter_io_out_0_aw_ready;
  wire  AXI4Fragmenter_io_out_0_aw_valid;
  wire [3:0] AXI4Fragmenter_io_out_0_aw_bits_id;
  wire [11:0] AXI4Fragmenter_io_out_0_aw_bits_addr;
  wire  AXI4Fragmenter_io_out_0_aw_bits_user;
  wire  AXI4Fragmenter_io_out_0_w_ready;
  wire  AXI4Fragmenter_io_out_0_w_valid;
  wire [63:0] AXI4Fragmenter_io_out_0_w_bits_data;
  wire [7:0] AXI4Fragmenter_io_out_0_w_bits_strb;
  wire  AXI4Fragmenter_io_out_0_w_bits_last;
  wire  AXI4Fragmenter_io_out_0_b_ready;
  wire  AXI4Fragmenter_io_out_0_b_valid;
  wire [3:0] AXI4Fragmenter_io_out_0_b_bits_id;
  wire [1:0] AXI4Fragmenter_io_out_0_b_bits_resp;
  wire  AXI4Fragmenter_io_out_0_b_bits_user;
  wire  AXI4Fragmenter_io_out_0_ar_ready;
  wire  AXI4Fragmenter_io_out_0_ar_valid;
  wire [3:0] AXI4Fragmenter_io_out_0_ar_bits_id;
  wire [11:0] AXI4Fragmenter_io_out_0_ar_bits_addr;
  wire  AXI4Fragmenter_io_out_0_ar_bits_user;
  wire  AXI4Fragmenter_io_out_0_r_ready;
  wire  AXI4Fragmenter_io_out_0_r_valid;
  wire [3:0] AXI4Fragmenter_io_out_0_r_bits_id;
  wire [63:0] AXI4Fragmenter_io_out_0_r_bits_data;
  wire [1:0] AXI4Fragmenter_io_out_0_r_bits_resp;
  wire  AXI4Fragmenter_io_out_0_r_bits_user;
  wire  AXI4Fragmenter_io_out_0_r_bits_last;
  wire  AXI4Buffer_clock;
  wire  AXI4Buffer_reset;
  wire  AXI4Buffer_io_in_0_aw_ready;
  wire  AXI4Buffer_io_in_0_aw_valid;
  wire [3:0] AXI4Buffer_io_in_0_aw_bits_id;
  wire [11:0] AXI4Buffer_io_in_0_aw_bits_addr;
  wire  AXI4Buffer_io_in_0_aw_bits_user;
  wire  AXI4Buffer_io_in_0_w_ready;
  wire  AXI4Buffer_io_in_0_w_valid;
  wire [63:0] AXI4Buffer_io_in_0_w_bits_data;
  wire [7:0] AXI4Buffer_io_in_0_w_bits_strb;
  wire  AXI4Buffer_io_in_0_w_bits_last;
  wire  AXI4Buffer_io_in_0_b_ready;
  wire  AXI4Buffer_io_in_0_b_valid;
  wire [3:0] AXI4Buffer_io_in_0_b_bits_id;
  wire [1:0] AXI4Buffer_io_in_0_b_bits_resp;
  wire  AXI4Buffer_io_in_0_b_bits_user;
  wire  AXI4Buffer_io_in_0_ar_ready;
  wire  AXI4Buffer_io_in_0_ar_valid;
  wire [3:0] AXI4Buffer_io_in_0_ar_bits_id;
  wire [11:0] AXI4Buffer_io_in_0_ar_bits_addr;
  wire  AXI4Buffer_io_in_0_ar_bits_user;
  wire  AXI4Buffer_io_in_0_r_ready;
  wire  AXI4Buffer_io_in_0_r_valid;
  wire [3:0] AXI4Buffer_io_in_0_r_bits_id;
  wire [63:0] AXI4Buffer_io_in_0_r_bits_data;
  wire [1:0] AXI4Buffer_io_in_0_r_bits_resp;
  wire  AXI4Buffer_io_in_0_r_bits_user;
  wire  AXI4Buffer_io_in_0_r_bits_last;
  wire  AXI4Buffer_io_out_0_aw_ready;
  wire  AXI4Buffer_io_out_0_aw_valid;
  wire [3:0] AXI4Buffer_io_out_0_aw_bits_id;
  wire [11:0] AXI4Buffer_io_out_0_aw_bits_addr;
  wire  AXI4Buffer_io_out_0_aw_bits_user;
  wire  AXI4Buffer_io_out_0_w_ready;
  wire  AXI4Buffer_io_out_0_w_valid;
  wire [63:0] AXI4Buffer_io_out_0_w_bits_data;
  wire [7:0] AXI4Buffer_io_out_0_w_bits_strb;
  wire  AXI4Buffer_io_out_0_b_ready;
  wire  AXI4Buffer_io_out_0_b_valid;
  wire [3:0] AXI4Buffer_io_out_0_b_bits_id;
  wire [1:0] AXI4Buffer_io_out_0_b_bits_resp;
  wire  AXI4Buffer_io_out_0_b_bits_user;
  wire  AXI4Buffer_io_out_0_ar_ready;
  wire  AXI4Buffer_io_out_0_ar_valid;
  wire [3:0] AXI4Buffer_io_out_0_ar_bits_id;
  wire [11:0] AXI4Buffer_io_out_0_ar_bits_addr;
  wire  AXI4Buffer_io_out_0_ar_bits_user;
  wire  AXI4Buffer_io_out_0_r_ready;
  wire  AXI4Buffer_io_out_0_r_valid;
  wire [3:0] AXI4Buffer_io_out_0_r_bits_id;
  wire [63:0] AXI4Buffer_io_out_0_r_bits_data;
  wire [1:0] AXI4Buffer_io_out_0_r_bits_resp;
  wire  AXI4Buffer_io_out_0_r_bits_user;
  wire  AXI4Buffer_io_out_0_r_bits_last;
  AXI4RAM AXI4RAM (
    .clock(AXI4RAM_clock),
    .reset(AXI4RAM_reset),
    .io_in_0_aw_ready(AXI4RAM_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4RAM_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4RAM_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4RAM_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_user(AXI4RAM_io_in_0_aw_bits_user),
    .io_in_0_w_ready(AXI4RAM_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4RAM_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4RAM_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4RAM_io_in_0_w_bits_strb),
    .io_in_0_b_ready(AXI4RAM_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4RAM_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4RAM_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4RAM_io_in_0_b_bits_resp),
    .io_in_0_b_bits_user(AXI4RAM_io_in_0_b_bits_user),
    .io_in_0_ar_ready(AXI4RAM_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4RAM_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4RAM_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4RAM_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_user(AXI4RAM_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4RAM_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4RAM_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4RAM_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4RAM_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4RAM_io_in_0_r_bits_resp),
    .io_in_0_r_bits_user(AXI4RAM_io_in_0_r_bits_user),
    .io_in_0_r_bits_last(AXI4RAM_io_in_0_r_bits_last)
  );
  AXI4Fragmenter_1 AXI4Fragmenter (
    .clock(AXI4Fragmenter_clock),
    .reset(AXI4Fragmenter_reset),
    .io_in_0_aw_ready(AXI4Fragmenter_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4Fragmenter_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4Fragmenter_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4Fragmenter_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_len(AXI4Fragmenter_io_in_0_aw_bits_len),
    .io_in_0_aw_bits_size(AXI4Fragmenter_io_in_0_aw_bits_size),
    .io_in_0_aw_bits_burst(AXI4Fragmenter_io_in_0_aw_bits_burst),
    .io_in_0_w_ready(AXI4Fragmenter_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4Fragmenter_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4Fragmenter_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4Fragmenter_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4Fragmenter_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4Fragmenter_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4Fragmenter_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4Fragmenter_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4Fragmenter_io_in_0_b_bits_resp),
    .io_in_0_ar_ready(AXI4Fragmenter_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4Fragmenter_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4Fragmenter_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4Fragmenter_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_len(AXI4Fragmenter_io_in_0_ar_bits_len),
    .io_in_0_ar_bits_size(AXI4Fragmenter_io_in_0_ar_bits_size),
    .io_in_0_ar_bits_burst(AXI4Fragmenter_io_in_0_ar_bits_burst),
    .io_in_0_r_ready(AXI4Fragmenter_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4Fragmenter_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4Fragmenter_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4Fragmenter_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4Fragmenter_io_in_0_r_bits_resp),
    .io_in_0_r_bits_last(AXI4Fragmenter_io_in_0_r_bits_last),
    .io_out_0_aw_ready(AXI4Fragmenter_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4Fragmenter_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4Fragmenter_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4Fragmenter_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_user(AXI4Fragmenter_io_out_0_aw_bits_user),
    .io_out_0_w_ready(AXI4Fragmenter_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4Fragmenter_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4Fragmenter_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4Fragmenter_io_out_0_w_bits_strb),
    .io_out_0_w_bits_last(AXI4Fragmenter_io_out_0_w_bits_last),
    .io_out_0_b_ready(AXI4Fragmenter_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4Fragmenter_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4Fragmenter_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(AXI4Fragmenter_io_out_0_b_bits_resp),
    .io_out_0_b_bits_user(AXI4Fragmenter_io_out_0_b_bits_user),
    .io_out_0_ar_ready(AXI4Fragmenter_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4Fragmenter_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4Fragmenter_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4Fragmenter_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_user(AXI4Fragmenter_io_out_0_ar_bits_user),
    .io_out_0_r_ready(AXI4Fragmenter_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4Fragmenter_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4Fragmenter_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(AXI4Fragmenter_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(AXI4Fragmenter_io_out_0_r_bits_resp),
    .io_out_0_r_bits_user(AXI4Fragmenter_io_out_0_r_bits_user),
    .io_out_0_r_bits_last(AXI4Fragmenter_io_out_0_r_bits_last)
  );
  AXI4Buffer_1 AXI4Buffer (
    .clock(AXI4Buffer_clock),
    .reset(AXI4Buffer_reset),
    .io_in_0_aw_ready(AXI4Buffer_io_in_0_aw_ready),
    .io_in_0_aw_valid(AXI4Buffer_io_in_0_aw_valid),
    .io_in_0_aw_bits_id(AXI4Buffer_io_in_0_aw_bits_id),
    .io_in_0_aw_bits_addr(AXI4Buffer_io_in_0_aw_bits_addr),
    .io_in_0_aw_bits_user(AXI4Buffer_io_in_0_aw_bits_user),
    .io_in_0_w_ready(AXI4Buffer_io_in_0_w_ready),
    .io_in_0_w_valid(AXI4Buffer_io_in_0_w_valid),
    .io_in_0_w_bits_data(AXI4Buffer_io_in_0_w_bits_data),
    .io_in_0_w_bits_strb(AXI4Buffer_io_in_0_w_bits_strb),
    .io_in_0_w_bits_last(AXI4Buffer_io_in_0_w_bits_last),
    .io_in_0_b_ready(AXI4Buffer_io_in_0_b_ready),
    .io_in_0_b_valid(AXI4Buffer_io_in_0_b_valid),
    .io_in_0_b_bits_id(AXI4Buffer_io_in_0_b_bits_id),
    .io_in_0_b_bits_resp(AXI4Buffer_io_in_0_b_bits_resp),
    .io_in_0_b_bits_user(AXI4Buffer_io_in_0_b_bits_user),
    .io_in_0_ar_ready(AXI4Buffer_io_in_0_ar_ready),
    .io_in_0_ar_valid(AXI4Buffer_io_in_0_ar_valid),
    .io_in_0_ar_bits_id(AXI4Buffer_io_in_0_ar_bits_id),
    .io_in_0_ar_bits_addr(AXI4Buffer_io_in_0_ar_bits_addr),
    .io_in_0_ar_bits_user(AXI4Buffer_io_in_0_ar_bits_user),
    .io_in_0_r_ready(AXI4Buffer_io_in_0_r_ready),
    .io_in_0_r_valid(AXI4Buffer_io_in_0_r_valid),
    .io_in_0_r_bits_id(AXI4Buffer_io_in_0_r_bits_id),
    .io_in_0_r_bits_data(AXI4Buffer_io_in_0_r_bits_data),
    .io_in_0_r_bits_resp(AXI4Buffer_io_in_0_r_bits_resp),
    .io_in_0_r_bits_user(AXI4Buffer_io_in_0_r_bits_user),
    .io_in_0_r_bits_last(AXI4Buffer_io_in_0_r_bits_last),
    .io_out_0_aw_ready(AXI4Buffer_io_out_0_aw_ready),
    .io_out_0_aw_valid(AXI4Buffer_io_out_0_aw_valid),
    .io_out_0_aw_bits_id(AXI4Buffer_io_out_0_aw_bits_id),
    .io_out_0_aw_bits_addr(AXI4Buffer_io_out_0_aw_bits_addr),
    .io_out_0_aw_bits_user(AXI4Buffer_io_out_0_aw_bits_user),
    .io_out_0_w_ready(AXI4Buffer_io_out_0_w_ready),
    .io_out_0_w_valid(AXI4Buffer_io_out_0_w_valid),
    .io_out_0_w_bits_data(AXI4Buffer_io_out_0_w_bits_data),
    .io_out_0_w_bits_strb(AXI4Buffer_io_out_0_w_bits_strb),
    .io_out_0_b_ready(AXI4Buffer_io_out_0_b_ready),
    .io_out_0_b_valid(AXI4Buffer_io_out_0_b_valid),
    .io_out_0_b_bits_id(AXI4Buffer_io_out_0_b_bits_id),
    .io_out_0_b_bits_resp(AXI4Buffer_io_out_0_b_bits_resp),
    .io_out_0_b_bits_user(AXI4Buffer_io_out_0_b_bits_user),
    .io_out_0_ar_ready(AXI4Buffer_io_out_0_ar_ready),
    .io_out_0_ar_valid(AXI4Buffer_io_out_0_ar_valid),
    .io_out_0_ar_bits_id(AXI4Buffer_io_out_0_ar_bits_id),
    .io_out_0_ar_bits_addr(AXI4Buffer_io_out_0_ar_bits_addr),
    .io_out_0_ar_bits_user(AXI4Buffer_io_out_0_ar_bits_user),
    .io_out_0_r_ready(AXI4Buffer_io_out_0_r_ready),
    .io_out_0_r_valid(AXI4Buffer_io_out_0_r_valid),
    .io_out_0_r_bits_id(AXI4Buffer_io_out_0_r_bits_id),
    .io_out_0_r_bits_data(AXI4Buffer_io_out_0_r_bits_data),
    .io_out_0_r_bits_resp(AXI4Buffer_io_out_0_r_bits_resp),
    .io_out_0_r_bits_user(AXI4Buffer_io_out_0_r_bits_user),
    .io_out_0_r_bits_last(AXI4Buffer_io_out_0_r_bits_last)
  );
  assign io_axi4_0_aw_ready = AXI4Fragmenter_io_in_0_aw_ready;
  assign io_axi4_0_w_ready = AXI4Fragmenter_io_in_0_w_ready;
  assign io_axi4_0_b_valid = AXI4Fragmenter_io_in_0_b_valid;
  assign io_axi4_0_b_bits_id = AXI4Fragmenter_io_in_0_b_bits_id;
  assign io_axi4_0_b_bits_resp = AXI4Fragmenter_io_in_0_b_bits_resp;
  assign io_axi4_0_ar_ready = AXI4Fragmenter_io_in_0_ar_ready;
  assign io_axi4_0_r_valid = AXI4Fragmenter_io_in_0_r_valid;
  assign io_axi4_0_r_bits_id = AXI4Fragmenter_io_in_0_r_bits_id;
  assign io_axi4_0_r_bits_data = AXI4Fragmenter_io_in_0_r_bits_data;
  assign io_axi4_0_r_bits_resp = AXI4Fragmenter_io_in_0_r_bits_resp;
  assign io_axi4_0_r_bits_last = AXI4Fragmenter_io_in_0_r_bits_last;
  assign AXI4RAM_clock = clock;
  assign AXI4RAM_reset = reset;
  assign AXI4RAM_io_in_0_aw_valid = AXI4Buffer_io_out_0_aw_valid;
  assign AXI4RAM_io_in_0_aw_bits_id = AXI4Buffer_io_out_0_aw_bits_id;
  assign AXI4RAM_io_in_0_aw_bits_addr = AXI4Buffer_io_out_0_aw_bits_addr;
  assign AXI4RAM_io_in_0_aw_bits_user = AXI4Buffer_io_out_0_aw_bits_user;
  assign AXI4RAM_io_in_0_w_valid = AXI4Buffer_io_out_0_w_valid;
  assign AXI4RAM_io_in_0_w_bits_data = AXI4Buffer_io_out_0_w_bits_data;
  assign AXI4RAM_io_in_0_w_bits_strb = AXI4Buffer_io_out_0_w_bits_strb;
  assign AXI4RAM_io_in_0_b_ready = AXI4Buffer_io_out_0_b_ready;
  assign AXI4RAM_io_in_0_ar_valid = AXI4Buffer_io_out_0_ar_valid;
  assign AXI4RAM_io_in_0_ar_bits_id = AXI4Buffer_io_out_0_ar_bits_id;
  assign AXI4RAM_io_in_0_ar_bits_addr = AXI4Buffer_io_out_0_ar_bits_addr;
  assign AXI4RAM_io_in_0_ar_bits_user = AXI4Buffer_io_out_0_ar_bits_user;
  assign AXI4RAM_io_in_0_r_ready = AXI4Buffer_io_out_0_r_ready;
  assign AXI4Fragmenter_clock = clock;
  assign AXI4Fragmenter_reset = reset;
  assign AXI4Fragmenter_io_in_0_aw_valid = io_axi4_0_aw_valid;
  assign AXI4Fragmenter_io_in_0_aw_bits_id = io_axi4_0_aw_bits_id;
  assign AXI4Fragmenter_io_in_0_aw_bits_addr = io_axi4_0_aw_bits_addr;
  assign AXI4Fragmenter_io_in_0_aw_bits_len = io_axi4_0_aw_bits_len;
  assign AXI4Fragmenter_io_in_0_aw_bits_size = io_axi4_0_aw_bits_size;
  assign AXI4Fragmenter_io_in_0_aw_bits_burst = io_axi4_0_aw_bits_burst;
  assign AXI4Fragmenter_io_in_0_w_valid = io_axi4_0_w_valid;
  assign AXI4Fragmenter_io_in_0_w_bits_data = io_axi4_0_w_bits_data;
  assign AXI4Fragmenter_io_in_0_w_bits_strb = io_axi4_0_w_bits_strb;
  assign AXI4Fragmenter_io_in_0_w_bits_last = io_axi4_0_w_bits_last;
  assign AXI4Fragmenter_io_in_0_b_ready = io_axi4_0_b_ready;
  assign AXI4Fragmenter_io_in_0_ar_valid = io_axi4_0_ar_valid;
  assign AXI4Fragmenter_io_in_0_ar_bits_id = io_axi4_0_ar_bits_id;
  assign AXI4Fragmenter_io_in_0_ar_bits_addr = io_axi4_0_ar_bits_addr;
  assign AXI4Fragmenter_io_in_0_ar_bits_len = io_axi4_0_ar_bits_len;
  assign AXI4Fragmenter_io_in_0_ar_bits_size = io_axi4_0_ar_bits_size;
  assign AXI4Fragmenter_io_in_0_ar_bits_burst = io_axi4_0_ar_bits_burst;
  assign AXI4Fragmenter_io_in_0_r_ready = io_axi4_0_r_ready;
  assign AXI4Fragmenter_io_out_0_aw_ready = AXI4Buffer_io_in_0_aw_ready;
  assign AXI4Fragmenter_io_out_0_w_ready = AXI4Buffer_io_in_0_w_ready;
  assign AXI4Fragmenter_io_out_0_b_valid = AXI4Buffer_io_in_0_b_valid;
  assign AXI4Fragmenter_io_out_0_b_bits_id = AXI4Buffer_io_in_0_b_bits_id;
  assign AXI4Fragmenter_io_out_0_b_bits_resp = AXI4Buffer_io_in_0_b_bits_resp;
  assign AXI4Fragmenter_io_out_0_b_bits_user = AXI4Buffer_io_in_0_b_bits_user;
  assign AXI4Fragmenter_io_out_0_ar_ready = AXI4Buffer_io_in_0_ar_ready;
  assign AXI4Fragmenter_io_out_0_r_valid = AXI4Buffer_io_in_0_r_valid;
  assign AXI4Fragmenter_io_out_0_r_bits_id = AXI4Buffer_io_in_0_r_bits_id;
  assign AXI4Fragmenter_io_out_0_r_bits_data = AXI4Buffer_io_in_0_r_bits_data;
  assign AXI4Fragmenter_io_out_0_r_bits_resp = AXI4Buffer_io_in_0_r_bits_resp;
  assign AXI4Fragmenter_io_out_0_r_bits_user = AXI4Buffer_io_in_0_r_bits_user;
  assign AXI4Fragmenter_io_out_0_r_bits_last = AXI4Buffer_io_in_0_r_bits_last;
  assign AXI4Buffer_clock = clock;
  assign AXI4Buffer_reset = reset;
  assign AXI4Buffer_io_in_0_aw_valid = AXI4Fragmenter_io_out_0_aw_valid;
  assign AXI4Buffer_io_in_0_aw_bits_id = AXI4Fragmenter_io_out_0_aw_bits_id;
  assign AXI4Buffer_io_in_0_aw_bits_addr = AXI4Fragmenter_io_out_0_aw_bits_addr;
  assign AXI4Buffer_io_in_0_aw_bits_user = AXI4Fragmenter_io_out_0_aw_bits_user;
  assign AXI4Buffer_io_in_0_w_valid = AXI4Fragmenter_io_out_0_w_valid;
  assign AXI4Buffer_io_in_0_w_bits_data = AXI4Fragmenter_io_out_0_w_bits_data;
  assign AXI4Buffer_io_in_0_w_bits_strb = AXI4Fragmenter_io_out_0_w_bits_strb;
  assign AXI4Buffer_io_in_0_w_bits_last = AXI4Fragmenter_io_out_0_w_bits_last;
  assign AXI4Buffer_io_in_0_b_ready = AXI4Fragmenter_io_out_0_b_ready;
  assign AXI4Buffer_io_in_0_ar_valid = AXI4Fragmenter_io_out_0_ar_valid;
  assign AXI4Buffer_io_in_0_ar_bits_id = AXI4Fragmenter_io_out_0_ar_bits_id;
  assign AXI4Buffer_io_in_0_ar_bits_addr = AXI4Fragmenter_io_out_0_ar_bits_addr;
  assign AXI4Buffer_io_in_0_ar_bits_user = AXI4Fragmenter_io_out_0_ar_bits_user;
  assign AXI4Buffer_io_in_0_r_ready = AXI4Fragmenter_io_out_0_r_ready;
  assign AXI4Buffer_io_out_0_aw_ready = AXI4RAM_io_in_0_aw_ready;
  assign AXI4Buffer_io_out_0_w_ready = AXI4RAM_io_in_0_w_ready;
  assign AXI4Buffer_io_out_0_b_valid = AXI4RAM_io_in_0_b_valid;
  assign AXI4Buffer_io_out_0_b_bits_id = AXI4RAM_io_in_0_b_bits_id;
  assign AXI4Buffer_io_out_0_b_bits_resp = AXI4RAM_io_in_0_b_bits_resp;
  assign AXI4Buffer_io_out_0_b_bits_user = AXI4RAM_io_in_0_b_bits_user;
  assign AXI4Buffer_io_out_0_ar_ready = AXI4RAM_io_in_0_ar_ready;
  assign AXI4Buffer_io_out_0_r_valid = AXI4RAM_io_in_0_r_valid;
  assign AXI4Buffer_io_out_0_r_bits_id = AXI4RAM_io_in_0_r_bits_id;
  assign AXI4Buffer_io_out_0_r_bits_data = AXI4RAM_io_in_0_r_bits_data;
  assign AXI4Buffer_io_out_0_r_bits_resp = AXI4RAM_io_in_0_r_bits_resp;
  assign AXI4Buffer_io_out_0_r_bits_user = AXI4RAM_io_in_0_r_bits_user;
  assign AXI4Buffer_io_out_0_r_bits_last = AXI4RAM_io_in_0_r_bits_last;
endmodule
module TestHarness(
  input   clock,
  input   reset,
  output  io_success
);
  wire  ExampleRocketSystem_clock;
  wire  ExampleRocketSystem_reset;
  wire  ExampleRocketSystem_debug_clockeddmi_dmi_req_ready;
  wire  ExampleRocketSystem_debug_clockeddmi_dmi_req_valid;
  wire [6:0] ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_addr;
  wire [31:0] ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_data;
  wire [1:0] ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_op;
  wire  ExampleRocketSystem_debug_clockeddmi_dmi_resp_ready;
  wire  ExampleRocketSystem_debug_clockeddmi_dmi_resp_valid;
  wire [31:0] ExampleRocketSystem_debug_clockeddmi_dmi_resp_bits_data;
  wire [1:0] ExampleRocketSystem_debug_clockeddmi_dmi_resp_bits_resp;
  wire  ExampleRocketSystem_debug_clockeddmi_dmiClock;
  wire  ExampleRocketSystem_debug_clockeddmi_dmiReset;
  wire  ExampleRocketSystem_debug_ndreset;
  wire [1:0] ExampleRocketSystem_interrupts;
  wire  ExampleRocketSystem_mmio_axi4_0_aw_ready;
  wire  ExampleRocketSystem_mmio_axi4_0_aw_valid;
  wire [3:0] ExampleRocketSystem_mmio_axi4_0_aw_bits_id;
  wire [30:0] ExampleRocketSystem_mmio_axi4_0_aw_bits_addr;
  wire [7:0] ExampleRocketSystem_mmio_axi4_0_aw_bits_len;
  wire [2:0] ExampleRocketSystem_mmio_axi4_0_aw_bits_size;
  wire [1:0] ExampleRocketSystem_mmio_axi4_0_aw_bits_burst;
  wire  ExampleRocketSystem_mmio_axi4_0_w_ready;
  wire  ExampleRocketSystem_mmio_axi4_0_w_valid;
  wire [63:0] ExampleRocketSystem_mmio_axi4_0_w_bits_data;
  wire [7:0] ExampleRocketSystem_mmio_axi4_0_w_bits_strb;
  wire  ExampleRocketSystem_mmio_axi4_0_w_bits_last;
  wire  ExampleRocketSystem_mmio_axi4_0_b_ready;
  wire  ExampleRocketSystem_mmio_axi4_0_b_valid;
  wire [3:0] ExampleRocketSystem_mmio_axi4_0_b_bits_id;
  wire [1:0] ExampleRocketSystem_mmio_axi4_0_b_bits_resp;
  wire  ExampleRocketSystem_mmio_axi4_0_ar_ready;
  wire  ExampleRocketSystem_mmio_axi4_0_ar_valid;
  wire [3:0] ExampleRocketSystem_mmio_axi4_0_ar_bits_id;
  wire [30:0] ExampleRocketSystem_mmio_axi4_0_ar_bits_addr;
  wire [7:0] ExampleRocketSystem_mmio_axi4_0_ar_bits_len;
  wire [2:0] ExampleRocketSystem_mmio_axi4_0_ar_bits_size;
  wire [1:0] ExampleRocketSystem_mmio_axi4_0_ar_bits_burst;
  wire  ExampleRocketSystem_mmio_axi4_0_r_ready;
  wire  ExampleRocketSystem_mmio_axi4_0_r_valid;
  wire [3:0] ExampleRocketSystem_mmio_axi4_0_r_bits_id;
  wire [63:0] ExampleRocketSystem_mmio_axi4_0_r_bits_data;
  wire [1:0] ExampleRocketSystem_mmio_axi4_0_r_bits_resp;
  wire  ExampleRocketSystem_mmio_axi4_0_r_bits_last;
  wire  ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_valid;
  wire [7:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_id;
  wire [31:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_addr;
  wire [7:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_len;
  wire [2:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_size;
  wire [1:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_burst;
  wire  ExampleRocketSystem_l2_frontend_bus_axi4_0_w_valid;
  wire [63:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_data;
  wire [7:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_strb;
  wire  ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_last;
  wire  ExampleRocketSystem_l2_frontend_bus_axi4_0_b_ready;
  wire  ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_valid;
  wire [7:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_id;
  wire [31:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_addr;
  wire [7:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_len;
  wire [2:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_size;
  wire [1:0] ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_burst;
  wire  ExampleRocketSystem_l2_frontend_bus_axi4_0_r_ready;
  wire  _T_3;
  wire  SimAXIMem_clock;
  wire  SimAXIMem_reset;
  wire  SimAXIMem_io_axi4_0_aw_ready;
  wire  SimAXIMem_io_axi4_0_aw_valid;
  wire [3:0] SimAXIMem_io_axi4_0_aw_bits_id;
  wire [11:0] SimAXIMem_io_axi4_0_aw_bits_addr;
  wire [7:0] SimAXIMem_io_axi4_0_aw_bits_len;
  wire [2:0] SimAXIMem_io_axi4_0_aw_bits_size;
  wire [1:0] SimAXIMem_io_axi4_0_aw_bits_burst;
  wire  SimAXIMem_io_axi4_0_w_ready;
  wire  SimAXIMem_io_axi4_0_w_valid;
  wire [63:0] SimAXIMem_io_axi4_0_w_bits_data;
  wire [7:0] SimAXIMem_io_axi4_0_w_bits_strb;
  wire  SimAXIMem_io_axi4_0_w_bits_last;
  wire  SimAXIMem_io_axi4_0_b_ready;
  wire  SimAXIMem_io_axi4_0_b_valid;
  wire [3:0] SimAXIMem_io_axi4_0_b_bits_id;
  wire [1:0] SimAXIMem_io_axi4_0_b_bits_resp;
  wire  SimAXIMem_io_axi4_0_ar_ready;
  wire  SimAXIMem_io_axi4_0_ar_valid;
  wire [3:0] SimAXIMem_io_axi4_0_ar_bits_id;
  wire [11:0] SimAXIMem_io_axi4_0_ar_bits_addr;
  wire [7:0] SimAXIMem_io_axi4_0_ar_bits_len;
  wire [2:0] SimAXIMem_io_axi4_0_ar_bits_size;
  wire [1:0] SimAXIMem_io_axi4_0_ar_bits_burst;
  wire  SimAXIMem_io_axi4_0_r_ready;
  wire  SimAXIMem_io_axi4_0_r_valid;
  wire [3:0] SimAXIMem_io_axi4_0_r_bits_id;
  wire [63:0] SimAXIMem_io_axi4_0_r_bits_data;
  wire [1:0] SimAXIMem_io_axi4_0_r_bits_resp;
  wire  SimAXIMem_io_axi4_0_r_bits_last;
  wire [31:0] SimDTM_exit;
  wire  SimDTM_debug_req_ready;
  wire  SimDTM_debug_req_valid;
  wire [6:0] SimDTM_debug_req_bits_addr;
  wire [31:0] SimDTM_debug_req_bits_data;
  wire [1:0] SimDTM_debug_req_bits_op;
  wire  SimDTM_debug_resp_ready;
  wire  SimDTM_debug_resp_valid;
  wire [31:0] SimDTM_debug_resp_bits_data;
  wire [1:0] SimDTM_debug_resp_bits_resp;
  wire  SimDTM_reset;
  wire  SimDTM_clk;
  wire  _T_11;
  wire  _T_13;
  wire [31:0] _T_15;
  wire  _T_17;
  ExampleRocketSystem ExampleRocketSystem (
    .clock(ExampleRocketSystem_clock),
    .reset(ExampleRocketSystem_reset),
    .debug_clockeddmi_dmi_req_ready(ExampleRocketSystem_debug_clockeddmi_dmi_req_ready),
    .debug_clockeddmi_dmi_req_valid(ExampleRocketSystem_debug_clockeddmi_dmi_req_valid),
    .debug_clockeddmi_dmi_req_bits_addr(ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_addr),
    .debug_clockeddmi_dmi_req_bits_data(ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_data),
    .debug_clockeddmi_dmi_req_bits_op(ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_op),
    .debug_clockeddmi_dmi_resp_ready(ExampleRocketSystem_debug_clockeddmi_dmi_resp_ready),
    .debug_clockeddmi_dmi_resp_valid(ExampleRocketSystem_debug_clockeddmi_dmi_resp_valid),
    .debug_clockeddmi_dmi_resp_bits_data(ExampleRocketSystem_debug_clockeddmi_dmi_resp_bits_data),
    .debug_clockeddmi_dmi_resp_bits_resp(ExampleRocketSystem_debug_clockeddmi_dmi_resp_bits_resp),
    .debug_clockeddmi_dmiClock(ExampleRocketSystem_debug_clockeddmi_dmiClock),
    .debug_clockeddmi_dmiReset(ExampleRocketSystem_debug_clockeddmi_dmiReset),
    .debug_ndreset(ExampleRocketSystem_debug_ndreset),
    .interrupts(ExampleRocketSystem_interrupts),
    .mmio_axi4_0_aw_ready(ExampleRocketSystem_mmio_axi4_0_aw_ready),
    .mmio_axi4_0_aw_valid(ExampleRocketSystem_mmio_axi4_0_aw_valid),
    .mmio_axi4_0_aw_bits_id(ExampleRocketSystem_mmio_axi4_0_aw_bits_id),
    .mmio_axi4_0_aw_bits_addr(ExampleRocketSystem_mmio_axi4_0_aw_bits_addr),
    .mmio_axi4_0_aw_bits_len(ExampleRocketSystem_mmio_axi4_0_aw_bits_len),
    .mmio_axi4_0_aw_bits_size(ExampleRocketSystem_mmio_axi4_0_aw_bits_size),
    .mmio_axi4_0_aw_bits_burst(ExampleRocketSystem_mmio_axi4_0_aw_bits_burst),
    .mmio_axi4_0_w_ready(ExampleRocketSystem_mmio_axi4_0_w_ready),
    .mmio_axi4_0_w_valid(ExampleRocketSystem_mmio_axi4_0_w_valid),
    .mmio_axi4_0_w_bits_data(ExampleRocketSystem_mmio_axi4_0_w_bits_data),
    .mmio_axi4_0_w_bits_strb(ExampleRocketSystem_mmio_axi4_0_w_bits_strb),
    .mmio_axi4_0_w_bits_last(ExampleRocketSystem_mmio_axi4_0_w_bits_last),
    .mmio_axi4_0_b_ready(ExampleRocketSystem_mmio_axi4_0_b_ready),
    .mmio_axi4_0_b_valid(ExampleRocketSystem_mmio_axi4_0_b_valid),
    .mmio_axi4_0_b_bits_id(ExampleRocketSystem_mmio_axi4_0_b_bits_id),
    .mmio_axi4_0_b_bits_resp(ExampleRocketSystem_mmio_axi4_0_b_bits_resp),
    .mmio_axi4_0_ar_ready(ExampleRocketSystem_mmio_axi4_0_ar_ready),
    .mmio_axi4_0_ar_valid(ExampleRocketSystem_mmio_axi4_0_ar_valid),
    .mmio_axi4_0_ar_bits_id(ExampleRocketSystem_mmio_axi4_0_ar_bits_id),
    .mmio_axi4_0_ar_bits_addr(ExampleRocketSystem_mmio_axi4_0_ar_bits_addr),
    .mmio_axi4_0_ar_bits_len(ExampleRocketSystem_mmio_axi4_0_ar_bits_len),
    .mmio_axi4_0_ar_bits_size(ExampleRocketSystem_mmio_axi4_0_ar_bits_size),
    .mmio_axi4_0_ar_bits_burst(ExampleRocketSystem_mmio_axi4_0_ar_bits_burst),
    .mmio_axi4_0_r_ready(ExampleRocketSystem_mmio_axi4_0_r_ready),
    .mmio_axi4_0_r_valid(ExampleRocketSystem_mmio_axi4_0_r_valid),
    .mmio_axi4_0_r_bits_id(ExampleRocketSystem_mmio_axi4_0_r_bits_id),
    .mmio_axi4_0_r_bits_data(ExampleRocketSystem_mmio_axi4_0_r_bits_data),
    .mmio_axi4_0_r_bits_resp(ExampleRocketSystem_mmio_axi4_0_r_bits_resp),
    .mmio_axi4_0_r_bits_last(ExampleRocketSystem_mmio_axi4_0_r_bits_last),
    .l2_frontend_bus_axi4_0_aw_valid(ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_valid),
    .l2_frontend_bus_axi4_0_aw_bits_id(ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_id),
    .l2_frontend_bus_axi4_0_aw_bits_addr(ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_addr),
    .l2_frontend_bus_axi4_0_aw_bits_len(ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_len),
    .l2_frontend_bus_axi4_0_aw_bits_size(ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_size),
    .l2_frontend_bus_axi4_0_aw_bits_burst(ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_burst),
    .l2_frontend_bus_axi4_0_w_valid(ExampleRocketSystem_l2_frontend_bus_axi4_0_w_valid),
    .l2_frontend_bus_axi4_0_w_bits_data(ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_data),
    .l2_frontend_bus_axi4_0_w_bits_strb(ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_strb),
    .l2_frontend_bus_axi4_0_w_bits_last(ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_last),
    .l2_frontend_bus_axi4_0_b_ready(ExampleRocketSystem_l2_frontend_bus_axi4_0_b_ready),
    .l2_frontend_bus_axi4_0_ar_valid(ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_valid),
    .l2_frontend_bus_axi4_0_ar_bits_id(ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_id),
    .l2_frontend_bus_axi4_0_ar_bits_addr(ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_addr),
    .l2_frontend_bus_axi4_0_ar_bits_len(ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_len),
    .l2_frontend_bus_axi4_0_ar_bits_size(ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_size),
    .l2_frontend_bus_axi4_0_ar_bits_burst(ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_burst),
    .l2_frontend_bus_axi4_0_r_ready(ExampleRocketSystem_l2_frontend_bus_axi4_0_r_ready)
  );
  SimAXIMem SimAXIMem (
    .clock(SimAXIMem_clock),
    .reset(SimAXIMem_reset),
    .io_axi4_0_aw_ready(SimAXIMem_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid(SimAXIMem_io_axi4_0_aw_valid),
    .io_axi4_0_aw_bits_id(SimAXIMem_io_axi4_0_aw_bits_id),
    .io_axi4_0_aw_bits_addr(SimAXIMem_io_axi4_0_aw_bits_addr),
    .io_axi4_0_aw_bits_len(SimAXIMem_io_axi4_0_aw_bits_len),
    .io_axi4_0_aw_bits_size(SimAXIMem_io_axi4_0_aw_bits_size),
    .io_axi4_0_aw_bits_burst(SimAXIMem_io_axi4_0_aw_bits_burst),
    .io_axi4_0_w_ready(SimAXIMem_io_axi4_0_w_ready),
    .io_axi4_0_w_valid(SimAXIMem_io_axi4_0_w_valid),
    .io_axi4_0_w_bits_data(SimAXIMem_io_axi4_0_w_bits_data),
    .io_axi4_0_w_bits_strb(SimAXIMem_io_axi4_0_w_bits_strb),
    .io_axi4_0_w_bits_last(SimAXIMem_io_axi4_0_w_bits_last),
    .io_axi4_0_b_ready(SimAXIMem_io_axi4_0_b_ready),
    .io_axi4_0_b_valid(SimAXIMem_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id(SimAXIMem_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp(SimAXIMem_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready(SimAXIMem_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid(SimAXIMem_io_axi4_0_ar_valid),
    .io_axi4_0_ar_bits_id(SimAXIMem_io_axi4_0_ar_bits_id),
    .io_axi4_0_ar_bits_addr(SimAXIMem_io_axi4_0_ar_bits_addr),
    .io_axi4_0_ar_bits_len(SimAXIMem_io_axi4_0_ar_bits_len),
    .io_axi4_0_ar_bits_size(SimAXIMem_io_axi4_0_ar_bits_size),
    .io_axi4_0_ar_bits_burst(SimAXIMem_io_axi4_0_ar_bits_burst),
    .io_axi4_0_r_ready(SimAXIMem_io_axi4_0_r_ready),
    .io_axi4_0_r_valid(SimAXIMem_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id(SimAXIMem_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data(SimAXIMem_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp(SimAXIMem_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last(SimAXIMem_io_axi4_0_r_bits_last)
  );
  SimDTM SimDTM (
    .exit(SimDTM_exit),
    .debug_req_ready(SimDTM_debug_req_ready),
    .debug_req_valid(SimDTM_debug_req_valid),
    .debug_req_bits_addr(SimDTM_debug_req_bits_addr),
    .debug_req_bits_data(SimDTM_debug_req_bits_data),
    .debug_req_bits_op(SimDTM_debug_req_bits_op),
    .debug_resp_ready(SimDTM_debug_resp_ready),
    .debug_resp_valid(SimDTM_debug_resp_valid),
    .debug_resp_bits_data(SimDTM_debug_resp_bits_data),
    .debug_resp_bits_resp(SimDTM_debug_resp_bits_resp),
    .reset(SimDTM_reset),
    .clk(SimDTM_clk)
  );
  assign io_success = _T_11;
  assign ExampleRocketSystem_clock = clock;
  assign ExampleRocketSystem_reset = _T_3;
  assign ExampleRocketSystem_debug_clockeddmi_dmi_req_valid = SimDTM_debug_req_valid;
  assign ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_addr = SimDTM_debug_req_bits_addr;
  assign ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_data = SimDTM_debug_req_bits_data;
  assign ExampleRocketSystem_debug_clockeddmi_dmi_req_bits_op = SimDTM_debug_req_bits_op;
  assign ExampleRocketSystem_debug_clockeddmi_dmi_resp_ready = SimDTM_debug_resp_ready;
  assign ExampleRocketSystem_debug_clockeddmi_dmiClock = clock;
  assign ExampleRocketSystem_debug_clockeddmi_dmiReset = reset;
  assign ExampleRocketSystem_interrupts = 2'h0;
  assign ExampleRocketSystem_mmio_axi4_0_aw_ready = SimAXIMem_io_axi4_0_aw_ready;
  assign ExampleRocketSystem_mmio_axi4_0_w_ready = SimAXIMem_io_axi4_0_w_ready;
  assign ExampleRocketSystem_mmio_axi4_0_b_valid = SimAXIMem_io_axi4_0_b_valid;
  assign ExampleRocketSystem_mmio_axi4_0_b_bits_id = SimAXIMem_io_axi4_0_b_bits_id;
  assign ExampleRocketSystem_mmio_axi4_0_b_bits_resp = SimAXIMem_io_axi4_0_b_bits_resp;
  assign ExampleRocketSystem_mmio_axi4_0_ar_ready = SimAXIMem_io_axi4_0_ar_ready;
  assign ExampleRocketSystem_mmio_axi4_0_r_valid = SimAXIMem_io_axi4_0_r_valid;
  assign ExampleRocketSystem_mmio_axi4_0_r_bits_id = SimAXIMem_io_axi4_0_r_bits_id;
  assign ExampleRocketSystem_mmio_axi4_0_r_bits_data = SimAXIMem_io_axi4_0_r_bits_data;
  assign ExampleRocketSystem_mmio_axi4_0_r_bits_resp = SimAXIMem_io_axi4_0_r_bits_resp;
  assign ExampleRocketSystem_mmio_axi4_0_r_bits_last = SimAXIMem_io_axi4_0_r_bits_last;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_valid = 1'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_id = 8'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_addr = 32'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_len = 8'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_size = 3'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_aw_bits_burst = 2'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_w_valid = 1'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_data = 64'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_strb = 8'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_w_bits_last = 1'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_b_ready = 1'h1;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_valid = 1'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_id = 8'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_addr = 32'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_len = 8'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_size = 3'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_ar_bits_burst = 2'h0;
  assign ExampleRocketSystem_l2_frontend_bus_axi4_0_r_ready = 1'h1;
  assign _T_3 = reset | ExampleRocketSystem_debug_ndreset;
  assign SimAXIMem_clock = clock;
  assign SimAXIMem_reset = reset;
  assign SimAXIMem_io_axi4_0_aw_valid = ExampleRocketSystem_mmio_axi4_0_aw_valid;
  assign SimAXIMem_io_axi4_0_aw_bits_id = ExampleRocketSystem_mmio_axi4_0_aw_bits_id;
  assign SimAXIMem_io_axi4_0_aw_bits_addr = ExampleRocketSystem_mmio_axi4_0_aw_bits_addr[11:0];
  assign SimAXIMem_io_axi4_0_aw_bits_len = ExampleRocketSystem_mmio_axi4_0_aw_bits_len;
  assign SimAXIMem_io_axi4_0_aw_bits_size = ExampleRocketSystem_mmio_axi4_0_aw_bits_size;
  assign SimAXIMem_io_axi4_0_aw_bits_burst = ExampleRocketSystem_mmio_axi4_0_aw_bits_burst;
  assign SimAXIMem_io_axi4_0_w_valid = ExampleRocketSystem_mmio_axi4_0_w_valid;
  assign SimAXIMem_io_axi4_0_w_bits_data = ExampleRocketSystem_mmio_axi4_0_w_bits_data;
  assign SimAXIMem_io_axi4_0_w_bits_strb = ExampleRocketSystem_mmio_axi4_0_w_bits_strb;
  assign SimAXIMem_io_axi4_0_w_bits_last = ExampleRocketSystem_mmio_axi4_0_w_bits_last;
  assign SimAXIMem_io_axi4_0_b_ready = ExampleRocketSystem_mmio_axi4_0_b_ready;
  assign SimAXIMem_io_axi4_0_ar_valid = ExampleRocketSystem_mmio_axi4_0_ar_valid;
  assign SimAXIMem_io_axi4_0_ar_bits_id = ExampleRocketSystem_mmio_axi4_0_ar_bits_id;
  assign SimAXIMem_io_axi4_0_ar_bits_addr = ExampleRocketSystem_mmio_axi4_0_ar_bits_addr[11:0];
  assign SimAXIMem_io_axi4_0_ar_bits_len = ExampleRocketSystem_mmio_axi4_0_ar_bits_len;
  assign SimAXIMem_io_axi4_0_ar_bits_size = ExampleRocketSystem_mmio_axi4_0_ar_bits_size;
  assign SimAXIMem_io_axi4_0_ar_bits_burst = ExampleRocketSystem_mmio_axi4_0_ar_bits_burst;
  assign SimAXIMem_io_axi4_0_r_ready = ExampleRocketSystem_mmio_axi4_0_r_ready;
  assign SimDTM_debug_req_ready = ExampleRocketSystem_debug_clockeddmi_dmi_req_ready;
  assign SimDTM_debug_resp_valid = ExampleRocketSystem_debug_clockeddmi_dmi_resp_valid;
  assign SimDTM_debug_resp_bits_data = ExampleRocketSystem_debug_clockeddmi_dmi_resp_bits_data;
  assign SimDTM_debug_resp_bits_resp = ExampleRocketSystem_debug_clockeddmi_dmi_resp_bits_resp;
  assign SimDTM_reset = reset;
  assign SimDTM_clk = clock;
  assign _T_11 = SimDTM_exit == 32'h1;
  assign _T_13 = SimDTM_exit >= 32'h2;
  assign _T_15 = SimDTM_exit >> 1'h1;
  assign _T_17 = reset == 1'h0;
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & _T_17) begin
          $fwrite(32'h80000002,"*** FAILED *** (exit code = %d)\n",_T_15);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13 & _T_17) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module data_arrays_0(
  input  [11:0] RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [7:0]  RW0_wdata_0,
  input  [7:0]  RW0_wdata_1,
  input  [7:0]  RW0_wdata_2,
  input  [7:0]  RW0_wdata_3,
  output [7:0]  RW0_rdata_0,
  output [7:0]  RW0_rdata_1,
  output [7:0]  RW0_rdata_2,
  output [7:0]  RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [11:0] data_arrays_0_ext_RW0_addr;
  wire  data_arrays_0_ext_RW0_en;
  wire  data_arrays_0_ext_RW0_clk;
  wire  data_arrays_0_ext_RW0_wmode;
  wire [31:0] data_arrays_0_ext_RW0_wdata;
  wire [31:0] data_arrays_0_ext_RW0_rdata;
  wire [3:0] data_arrays_0_ext_RW0_wmask;
  wire [7:0] _GEN_0;
  wire [7:0] _GEN_1;
  wire [7:0] _GEN_2;
  wire [7:0] _GEN_3;
  wire [7:0] _GEN_4;
  wire [7:0] _GEN_5;
  wire [7:0] _GEN_6;
  wire [7:0] _GEN_7;
  wire [15:0] _GEN_8;
  wire [15:0] _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire [1:0] _GEN_14;
  wire [1:0] _GEN_15;
  data_arrays_0_ext data_arrays_0_ext (
    .RW0_addr(data_arrays_0_ext_RW0_addr),
    .RW0_en(data_arrays_0_ext_RW0_en),
    .RW0_clk(data_arrays_0_ext_RW0_clk),
    .RW0_wmode(data_arrays_0_ext_RW0_wmode),
    .RW0_wdata(data_arrays_0_ext_RW0_wdata),
    .RW0_rdata(data_arrays_0_ext_RW0_rdata),
    .RW0_wmask(data_arrays_0_ext_RW0_wmask)
  );
  assign RW0_rdata_0 = $unsigned(_GEN_0);
  assign RW0_rdata_1 = $unsigned(_GEN_1);
  assign RW0_rdata_2 = $unsigned(_GEN_2);
  assign RW0_rdata_3 = $unsigned(_GEN_3);
  assign data_arrays_0_ext_RW0_addr = RW0_addr;
  assign data_arrays_0_ext_RW0_en = RW0_en;
  assign data_arrays_0_ext_RW0_clk = RW0_clk;
  assign data_arrays_0_ext_RW0_wmode = RW0_wmode;
  assign data_arrays_0_ext_RW0_wdata = {_GEN_8,_GEN_9};
  assign data_arrays_0_ext_RW0_wmask = {_GEN_14,_GEN_15};
  assign _GEN_0 = data_arrays_0_ext_RW0_rdata[7:0];
  assign _GEN_1 = data_arrays_0_ext_RW0_rdata[15:8];
  assign _GEN_2 = data_arrays_0_ext_RW0_rdata[23:16];
  assign _GEN_3 = data_arrays_0_ext_RW0_rdata[31:24];
  assign _GEN_4 = $unsigned(RW0_wdata_3);
  assign _GEN_5 = $unsigned(RW0_wdata_2);
  assign _GEN_6 = $unsigned(RW0_wdata_1);
  assign _GEN_7 = $unsigned(RW0_wdata_0);
  assign _GEN_8 = {_GEN_4,_GEN_5};
  assign _GEN_9 = {_GEN_6,_GEN_7};
  assign _GEN_10 = $unsigned(RW0_wmask_3);
  assign _GEN_11 = $unsigned(RW0_wmask_2);
  assign _GEN_12 = $unsigned(RW0_wmask_1);
  assign _GEN_13 = $unsigned(RW0_wmask_0);
  assign _GEN_14 = {_GEN_10,_GEN_11};
  assign _GEN_15 = {_GEN_12,_GEN_13};
endmodule
module tag_array(
  input  [5:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [20:0] RW0_wdata_0,
  output [20:0] RW0_rdata_0,
  input         RW0_wmask_0
);
  wire [5:0] tag_array_ext_RW0_addr;
  wire  tag_array_ext_RW0_en;
  wire  tag_array_ext_RW0_clk;
  wire  tag_array_ext_RW0_wmode;
  wire [20:0] tag_array_ext_RW0_wdata;
  wire [20:0] tag_array_ext_RW0_rdata;
  wire  tag_array_ext_RW0_wmask;
  tag_array_ext tag_array_ext (
    .RW0_addr(tag_array_ext_RW0_addr),
    .RW0_en(tag_array_ext_RW0_en),
    .RW0_clk(tag_array_ext_RW0_clk),
    .RW0_wmode(tag_array_ext_RW0_wmode),
    .RW0_wdata(tag_array_ext_RW0_wdata),
    .RW0_rdata(tag_array_ext_RW0_rdata),
    .RW0_wmask(tag_array_ext_RW0_wmask)
  );
  assign RW0_rdata_0 = $unsigned(tag_array_ext_RW0_rdata);
  assign tag_array_ext_RW0_addr = RW0_addr;
  assign tag_array_ext_RW0_en = RW0_en;
  assign tag_array_ext_RW0_clk = RW0_clk;
  assign tag_array_ext_RW0_wmode = RW0_wmode;
  assign tag_array_ext_RW0_wdata = $unsigned(RW0_wdata_0);
  assign tag_array_ext_RW0_wmask = $unsigned(RW0_wmask_0);
endmodule
module data_arrays_0_0(
  input  [9:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [31:0] RW0_wdata_0,
  output [31:0] RW0_rdata_0,
  input         RW0_wmask_0
);
  wire [9:0] data_arrays_0_0_ext_RW0_addr;
  wire  data_arrays_0_0_ext_RW0_en;
  wire  data_arrays_0_0_ext_RW0_clk;
  wire  data_arrays_0_0_ext_RW0_wmode;
  wire [31:0] data_arrays_0_0_ext_RW0_wdata;
  wire [31:0] data_arrays_0_0_ext_RW0_rdata;
  wire  data_arrays_0_0_ext_RW0_wmask;
  data_arrays_0_0_ext data_arrays_0_0_ext (
    .RW0_addr(data_arrays_0_0_ext_RW0_addr),
    .RW0_en(data_arrays_0_0_ext_RW0_en),
    .RW0_clk(data_arrays_0_0_ext_RW0_clk),
    .RW0_wmode(data_arrays_0_0_ext_RW0_wmode),
    .RW0_wdata(data_arrays_0_0_ext_RW0_wdata),
    .RW0_rdata(data_arrays_0_0_ext_RW0_rdata),
    .RW0_wmask(data_arrays_0_0_ext_RW0_wmask)
  );
  assign RW0_rdata_0 = $unsigned(data_arrays_0_0_ext_RW0_rdata);
  assign data_arrays_0_0_ext_RW0_addr = RW0_addr;
  assign data_arrays_0_0_ext_RW0_en = RW0_en;
  assign data_arrays_0_0_ext_RW0_clk = RW0_clk;
  assign data_arrays_0_0_ext_RW0_wmode = RW0_wmode;
  assign data_arrays_0_0_ext_RW0_wdata = $unsigned(RW0_wdata_0);
  assign data_arrays_0_0_ext_RW0_wmask = $unsigned(RW0_wmask_0);
endmodule
module mem(
  input  [8:0] R0_addr,
  input        R0_en,
  input        R0_clk,
  output [7:0] R0_data_0,
  output [7:0] R0_data_1,
  output [7:0] R0_data_2,
  output [7:0] R0_data_3,
  output [7:0] R0_data_4,
  output [7:0] R0_data_5,
  output [7:0] R0_data_6,
  output [7:0] R0_data_7,
  input  [8:0] W0_addr,
  input        W0_en,
  input        W0_clk,
  input  [7:0] W0_data_0,
  input  [7:0] W0_data_1,
  input  [7:0] W0_data_2,
  input  [7:0] W0_data_3,
  input  [7:0] W0_data_4,
  input  [7:0] W0_data_5,
  input  [7:0] W0_data_6,
  input  [7:0] W0_data_7,
  input        W0_mask_0,
  input        W0_mask_1,
  input        W0_mask_2,
  input        W0_mask_3,
  input        W0_mask_4,
  input        W0_mask_5,
  input        W0_mask_6,
  input        W0_mask_7
);
  wire [8:0] mem_ext_R0_addr;
  wire  mem_ext_R0_en;
  wire  mem_ext_R0_clk;
  wire [63:0] mem_ext_R0_data;
  wire [8:0] mem_ext_W0_addr;
  wire  mem_ext_W0_en;
  wire  mem_ext_W0_clk;
  wire [63:0] mem_ext_W0_data;
  wire [7:0] mem_ext_W0_mask;
  wire [7:0] _GEN_0;
  wire [7:0] _GEN_1;
  wire [7:0] _GEN_2;
  wire [7:0] _GEN_3;
  wire [7:0] _GEN_4;
  wire [7:0] _GEN_5;
  wire [7:0] _GEN_6;
  wire [7:0] _GEN_7;
  wire [7:0] _GEN_8;
  wire [7:0] _GEN_9;
  wire [7:0] _GEN_10;
  wire [7:0] _GEN_11;
  wire [15:0] _GEN_12;
  wire [15:0] _GEN_13;
  wire [7:0] _GEN_14;
  wire [7:0] _GEN_15;
  wire [7:0] _GEN_16;
  wire [7:0] _GEN_17;
  wire [15:0] _GEN_18;
  wire [15:0] _GEN_19;
  wire [31:0] _GEN_20;
  wire [31:0] _GEN_21;
  wire  _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire  _GEN_25;
  wire [1:0] _GEN_26;
  wire [1:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire  _GEN_30;
  wire  _GEN_31;
  wire [1:0] _GEN_32;
  wire [1:0] _GEN_33;
  wire [3:0] _GEN_34;
  wire [3:0] _GEN_35;
  mem_ext mem_ext (
    .R0_addr(mem_ext_R0_addr),
    .R0_en(mem_ext_R0_en),
    .R0_clk(mem_ext_R0_clk),
    .R0_data(mem_ext_R0_data),
    .W0_addr(mem_ext_W0_addr),
    .W0_en(mem_ext_W0_en),
    .W0_clk(mem_ext_W0_clk),
    .W0_data(mem_ext_W0_data),
    .W0_mask(mem_ext_W0_mask)
  );
  assign R0_data_0 = $unsigned(_GEN_0);
  assign R0_data_1 = $unsigned(_GEN_1);
  assign R0_data_2 = $unsigned(_GEN_2);
  assign R0_data_3 = $unsigned(_GEN_3);
  assign R0_data_4 = $unsigned(_GEN_4);
  assign R0_data_5 = $unsigned(_GEN_5);
  assign R0_data_6 = $unsigned(_GEN_6);
  assign R0_data_7 = $unsigned(_GEN_7);
  assign mem_ext_R0_addr = R0_addr;
  assign mem_ext_R0_en = R0_en;
  assign mem_ext_R0_clk = R0_clk;
  assign mem_ext_W0_addr = W0_addr;
  assign mem_ext_W0_en = W0_en;
  assign mem_ext_W0_clk = W0_clk;
  assign mem_ext_W0_data = {_GEN_20,_GEN_21};
  assign mem_ext_W0_mask = {_GEN_34,_GEN_35};
  assign _GEN_0 = mem_ext_R0_data[7:0];
  assign _GEN_1 = mem_ext_R0_data[15:8];
  assign _GEN_2 = mem_ext_R0_data[23:16];
  assign _GEN_3 = mem_ext_R0_data[31:24];
  assign _GEN_4 = mem_ext_R0_data[39:32];
  assign _GEN_5 = mem_ext_R0_data[47:40];
  assign _GEN_6 = mem_ext_R0_data[55:48];
  assign _GEN_7 = mem_ext_R0_data[63:56];
  assign _GEN_8 = $unsigned(W0_data_7);
  assign _GEN_9 = $unsigned(W0_data_6);
  assign _GEN_10 = $unsigned(W0_data_5);
  assign _GEN_11 = $unsigned(W0_data_4);
  assign _GEN_12 = {_GEN_8,_GEN_9};
  assign _GEN_13 = {_GEN_10,_GEN_11};
  assign _GEN_14 = $unsigned(W0_data_3);
  assign _GEN_15 = $unsigned(W0_data_2);
  assign _GEN_16 = $unsigned(W0_data_1);
  assign _GEN_17 = $unsigned(W0_data_0);
  assign _GEN_18 = {_GEN_14,_GEN_15};
  assign _GEN_19 = {_GEN_16,_GEN_17};
  assign _GEN_20 = {_GEN_12,_GEN_13};
  assign _GEN_21 = {_GEN_18,_GEN_19};
  assign _GEN_22 = $unsigned(W0_mask_7);
  assign _GEN_23 = $unsigned(W0_mask_6);
  assign _GEN_24 = $unsigned(W0_mask_5);
  assign _GEN_25 = $unsigned(W0_mask_4);
  assign _GEN_26 = {_GEN_22,_GEN_23};
  assign _GEN_27 = {_GEN_24,_GEN_25};
  assign _GEN_28 = $unsigned(W0_mask_3);
  assign _GEN_29 = $unsigned(W0_mask_2);
  assign _GEN_30 = $unsigned(W0_mask_1);
  assign _GEN_31 = $unsigned(W0_mask_0);
  assign _GEN_32 = {_GEN_28,_GEN_29};
  assign _GEN_33 = {_GEN_30,_GEN_31};
  assign _GEN_34 = {_GEN_26,_GEN_27};
  assign _GEN_35 = {_GEN_32,_GEN_33};
endmodule
